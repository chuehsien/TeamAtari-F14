module audioControl;


endmodule