module POKEYTest


endmodule