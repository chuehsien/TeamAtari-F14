module interruptControl


endmodule