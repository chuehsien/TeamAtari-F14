module interruptControlTest


endmodule