module randomLogic (T,OP,prevOP,phi1,phi2,activeInt,carry,statusC,decMode,control);
    input [6:0] T;
    input [7:0] OP,prevOP;
    input [2:0] activeInt;
    input phi1,phi2,carry,statusC,decMode;
    output [64:0] control;
    
    assign control[64:62] = 3'b000; //reserve for future use.
    
assign control[`DL_DB] = (OP==`BRK & T==`Tzero & phi1)
			 | (OP==`BRK & T==`Tzero & phi2)
			 | (OP==`BRK & T==`Tone & phi1)
			 | (OP==`BRK & T==`Tsix & phi2)
			 | (OP==`ORA_izx & T==`Tzero & phi2)
			 | (OP==`ORA_izx & T==`Tone & phi1)
			 | (OP==`ORA_izx & T==`Tthree & phi2)
			 | (OP==`ORA_izx & T==`Tfour & phi1)
			 | (OP==`ORA_izx & T==`Tfour & phi2)
			 | (OP==`ORA_izx & T==`Tfive & phi1)
			 | (OP==`ORA_zp & T==`Tzero & phi2)
			 | (OP==`ORA_zp & T==`Tone & phi1)
			 | (OP==`ASL_zp & T==`Tzero & phi2)
			 | (OP==`ASL_zp & T==`Tone & phi1)
			 | (OP==`ASL_zp & T==`Tthree & phi2)
			 | (OP==`ASL_zp & T==`Tfour & phi1)
			 | (OP==`PHP & T==`Tzero & phi2)
			 | (OP==`PHP & T==`Tone & phi1)
			 | (OP==`ORA_imm & T==`Tone & phi1)
			 | (OP==`ORA_imm & T==`Ttwo & phi2)
			 | (OP==`ORA_abs & T==`Tzero & phi2)
			 | (OP==`ORA_abs & T==`Tone & phi1)
			 | (OP==`ORA_abs & T==`Ttwo & phi2)
			 | (OP==`ORA_abs & T==`Tthree & phi1)
			 | (OP==`ASL_abs & T==`Tzero & phi2)
			 | (OP==`ASL_abs & T==`Tone & phi1)
			 | (OP==`ASL_abs & T==`Ttwo & phi2)
			 | (OP==`ASL_abs & T==`Tthree & phi1)
			 | (OP==`ASL_abs & T==`Tfour & phi2)
			 | (OP==`ASL_abs & T==`Tfive & phi1)
			 | (OP==`BPL_rel & T==`Tzero & phi2)
			 | (OP==`BPL_rel & T==`Ttwo & phi2)
			 | (OP==`BPL_rel & T==`Tthree & phi1)
			 | (OP==`BPL_rel & T==`T1BranchCross & phi1)
			 | (OP==`BPL_rel & T==`T1NoBranch & phi1)
			 | (OP==`ORA_izy & T==`TzeroCrossPg & phi2)
			 | (OP==`ORA_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ORA_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`ORA_izy & T==`Tone & phi1)
			 | (OP==`ORA_izy & T==`Ttwo & phi2)
			 | (OP==`ORA_izy & T==`Tthree & phi1)
			 | (OP==`ORA_izy & T==`Tthree & phi2)
			 | (OP==`ORA_izy & T==`Tfour & phi1)
			 | (OP==`ORA_izy & T==`Tfour & phi2)
			 | (OP==`ORA_izy & T==`Tfive & phi1)
			 | (OP==`ORA_zpx & T==`Tzero & phi2)
			 | (OP==`ORA_zpx & T==`Tone & phi1)
			 | (OP==`ASL_zpx & T==`Tzero & phi2)
			 | (OP==`ASL_zpx & T==`Tone & phi1)
			 | (OP==`ASL_zpx & T==`Tfour & phi2)
			 | (OP==`ASL_zpx & T==`Tfive & phi1)
			 | (OP==`ORA_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ORA_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`ORA_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`ORA_aby & T==`Tone & phi1)
			 | (OP==`ORA_aby & T==`Ttwo & phi2)
			 | (OP==`ORA_aby & T==`Tthree & phi1)
			 | (OP==`ORA_aby & T==`Tthree & phi2)
			 | (OP==`ORA_aby & T==`Tfour & phi1)
			 | (OP==`ORA_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ORA_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`ORA_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`ORA_abx & T==`Tone & phi1)
			 | (OP==`ORA_abx & T==`Ttwo & phi2)
			 | (OP==`ORA_abx & T==`Tthree & phi1)
			 | (OP==`ORA_abx & T==`Tthree & phi2)
			 | (OP==`ORA_abx & T==`Tfour & phi1)
			 | (OP==`ASL_abx & T==`Tzero & phi2)
			 | (OP==`ASL_abx & T==`Tone & phi1)
			 | (OP==`ASL_abx & T==`Ttwo & phi2)
			 | (OP==`ASL_abx & T==`Tthree & phi1)
			 | (OP==`ASL_abx & T==`Tthree & phi2)
			 | (OP==`ASL_abx & T==`Tfour & phi1)
			 | (OP==`ASL_abx & T==`Tfive & phi2)
			 | (OP==`ASL_abx & T==`Tsix & phi1)
			 | (OP==`JSR_abs & T==`Tzero & phi2)
			 | (OP==`JSR_abs & T==`Tone & phi1)
			 | (OP==`JSR_abs & T==`Ttwo & phi2)
			 | (OP==`JSR_abs & T==`Tthree & phi1)
			 | (OP==`AND_izx & T==`Tzero & phi2)
			 | (OP==`AND_izx & T==`Tone & phi1)
			 | (OP==`AND_izx & T==`Tthree & phi2)
			 | (OP==`AND_izx & T==`Tfour & phi1)
			 | (OP==`AND_izx & T==`Tfour & phi2)
			 | (OP==`AND_izx & T==`Tfive & phi1)
			 | (OP==`BIT_zp & T==`Tzero & phi2)
			 | (OP==`BIT_zp & T==`Tone & phi1)
			 | (OP==`AND_zp & T==`Tzero & phi2)
			 | (OP==`AND_zp & T==`Tone & phi1)
			 | (OP==`ROL_zp & T==`Tzero & phi2)
			 | (OP==`ROL_zp & T==`Tone & phi1)
			 | (OP==`ROL_zp & T==`Tthree & phi2)
			 | (OP==`ROL_zp & T==`Tfour & phi1)
			 | (OP==`PLP & T==`Tzero & phi1)
			 | (OP==`PLP & T==`Tzero & phi2)
			 | (OP==`PLP & T==`Tone & phi1)
			 | (OP==`PLP & T==`Tone & phi2)
			 | (OP==`PLP & T==`Ttwo & phi2)
			 | (OP==`PLP & T==`Tthree & phi1)
			 | (OP==`PLP & T==`Tthree & phi2)
			 | (OP==`AND_imm & T==`Tone & phi1)
			 | (OP==`AND_imm & T==`Ttwo & phi2)
			 | (OP==`BIT_abs & T==`Tzero & phi2)
			 | (OP==`BIT_abs & T==`Tone & phi1)
			 | (OP==`BIT_abs & T==`Ttwo & phi2)
			 | (OP==`BIT_abs & T==`Tthree & phi1)
			 | (OP==`AND_abs & T==`Tzero & phi2)
			 | (OP==`AND_abs & T==`Tone & phi1)
			 | (OP==`AND_abs & T==`Ttwo & phi2)
			 | (OP==`AND_abs & T==`Tthree & phi1)
			 | (OP==`ROL_abs & T==`Tzero & phi2)
			 | (OP==`ROL_abs & T==`Tone & phi1)
			 | (OP==`ROL_abs & T==`Ttwo & phi2)
			 | (OP==`ROL_abs & T==`Tthree & phi1)
			 | (OP==`ROL_abs & T==`Tfour & phi2)
			 | (OP==`ROL_abs & T==`Tfive & phi1)
			 | (OP==`BMI_rel & T==`Tzero & phi2)
			 | (OP==`BMI_rel & T==`Ttwo & phi2)
			 | (OP==`BMI_rel & T==`Tthree & phi1)
			 | (OP==`BMI_rel & T==`T1BranchCross & phi1)
			 | (OP==`BMI_rel & T==`T1NoBranch & phi1)
			 | (OP==`AND_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`AND_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`AND_izy & T==`TzeroCrossPg & phi2)
			 | (OP==`AND_izy & T==`Tone & phi1)
			 | (OP==`AND_izy & T==`Ttwo & phi2)
			 | (OP==`AND_izy & T==`Tthree & phi1)
			 | (OP==`AND_izy & T==`Tthree & phi2)
			 | (OP==`AND_izy & T==`Tfour & phi1)
			 | (OP==`AND_izy & T==`Tfour & phi2)
			 | (OP==`AND_izy & T==`Tfive & phi1)
			 | (OP==`AND_zpx & T==`Tzero & phi2)
			 | (OP==`AND_zpx & T==`Tone & phi1)
			 | (OP==`ROL_zpx & T==`Tzero & phi2)
			 | (OP==`ROL_zpx & T==`Tone & phi1)
			 | (OP==`ROL_zpx & T==`Tfour & phi2)
			 | (OP==`ROL_zpx & T==`Tfive & phi1)
			 | (OP==`AND_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`AND_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`AND_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`AND_aby & T==`Tone & phi1)
			 | (OP==`AND_aby & T==`Ttwo & phi2)
			 | (OP==`AND_aby & T==`Tthree & phi1)
			 | (OP==`AND_aby & T==`Tthree & phi2)
			 | (OP==`AND_aby & T==`Tfour & phi1)
			 | (OP==`AND_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`AND_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`AND_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`AND_abx & T==`Tone & phi1)
			 | (OP==`AND_abx & T==`Ttwo & phi2)
			 | (OP==`AND_abx & T==`Tthree & phi1)
			 | (OP==`AND_abx & T==`Tthree & phi2)
			 | (OP==`AND_abx & T==`Tfour & phi1)
			 | (OP==`ROL_abx & T==`Tzero & phi2)
			 | (OP==`ROL_abx & T==`Tone & phi1)
			 | (OP==`ROL_abx & T==`Ttwo & phi2)
			 | (OP==`ROL_abx & T==`Tthree & phi1)
			 | (OP==`ROL_abx & T==`Tthree & phi2)
			 | (OP==`ROL_abx & T==`Tfour & phi1)
			 | (OP==`ROL_abx & T==`Tfive & phi2)
			 | (OP==`ROL_abx & T==`Tsix & phi1)
			 | (OP==`RTI & T==`Tzero & phi1)
			 | (OP==`RTI & T==`Tzero & phi2)
			 | (OP==`RTI & T==`Tone & phi1)
			 | (OP==`RTI & T==`Tone & phi2)
			 | (OP==`RTI & T==`Ttwo & phi2)
			 | (OP==`RTI & T==`Tthree & phi1)
			 | (OP==`RTI & T==`Tthree & phi2)
			 | (OP==`RTI & T==`Tfour & phi1)
			 | (OP==`RTI & T==`Tfour & phi2)
			 | (OP==`RTI & T==`Tfive & phi1)
			 | (OP==`RTI & T==`Tfive & phi2)
			 | (OP==`EOR_izx & T==`Tzero & phi2)
			 | (OP==`EOR_izx & T==`Tone & phi1)
			 | (OP==`EOR_izx & T==`Tthree & phi2)
			 | (OP==`EOR_izx & T==`Tfour & phi1)
			 | (OP==`EOR_izx & T==`Tfour & phi2)
			 | (OP==`EOR_izx & T==`Tfive & phi1)
			 | (OP==`EOR_zp & T==`Tzero & phi2)
			 | (OP==`EOR_zp & T==`Tone & phi1)
			 | (OP==`LSR_zp & T==`Tzero & phi2)
			 | (OP==`LSR_zp & T==`Tone & phi1)
			 | (OP==`LSR_zp & T==`Tthree & phi2)
			 | (OP==`LSR_zp & T==`Tfour & phi1)
			 | (OP==`PHA & T==`Tzero & phi2)
			 | (OP==`PHA & T==`Tone & phi1)
			 | (OP==`EOR_imm & T==`Tone & phi1)
			 | (OP==`EOR_imm & T==`Ttwo & phi2)
			 | (OP==`JMP_abs & T==`Tzero & phi1)
			 | (OP==`JMP_abs & T==`Tzero & phi2)
			 | (OP==`JMP_abs & T==`Tone & phi1)
			 | (OP==`JMP_abs & T==`Ttwo & phi2)
			 | (OP==`EOR_abs & T==`Tzero & phi2)
			 | (OP==`EOR_abs & T==`Tone & phi1)
			 | (OP==`EOR_abs & T==`Ttwo & phi2)
			 | (OP==`EOR_abs & T==`Tthree & phi1)
			 | (OP==`LSR_abs & T==`Tzero & phi2)
			 | (OP==`LSR_abs & T==`Tone & phi1)
			 | (OP==`LSR_abs & T==`Ttwo & phi2)
			 | (OP==`LSR_abs & T==`Tthree & phi1)
			 | (OP==`LSR_abs & T==`Tfour & phi2)
			 | (OP==`LSR_abs & T==`Tfive & phi1)
			 | (OP==`BVC_rel & T==`Tzero & phi2)
			 | (OP==`BVC_rel & T==`Ttwo & phi2)
			 | (OP==`BVC_rel & T==`Tthree & phi1)
			 | (OP==`BVC_rel & T==`T1BranchCross & phi1)
			 | (OP==`BVC_rel & T==`T1NoBranch & phi1)
			 | (OP==`EOR_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`EOR_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`EOR_izy & T==`TzeroCrossPg & phi2)
			 | (OP==`EOR_izy & T==`Tone & phi1)
			 | (OP==`EOR_izy & T==`Ttwo & phi2)
			 | (OP==`EOR_izy & T==`Tthree & phi1)
			 | (OP==`EOR_izy & T==`Tthree & phi2)
			 | (OP==`EOR_izy & T==`Tfour & phi1)
			 | (OP==`EOR_izy & T==`Tfour & phi2)
			 | (OP==`EOR_izy & T==`Tfive & phi1)
			 | (OP==`EOR_zpx & T==`Tzero & phi2)
			 | (OP==`EOR_zpx & T==`Tone & phi1)
			 | (OP==`LSR_zpx & T==`Tzero & phi2)
			 | (OP==`LSR_zpx & T==`Tone & phi1)
			 | (OP==`LSR_zpx & T==`Tfour & phi2)
			 | (OP==`LSR_zpx & T==`Tfive & phi1)
			 | (OP==`EOR_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`EOR_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`EOR_aby & T==`Tone & phi1)
			 | (OP==`EOR_aby & T==`Ttwo & phi2)
			 | (OP==`EOR_aby & T==`Tthree & phi1)
			 | (OP==`EOR_aby & T==`Tthree & phi2)
			 | (OP==`EOR_aby & T==`Tfour & phi1)
			 | (OP==`EOR_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`EOR_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`EOR_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`EOR_abx & T==`Tone & phi1)
			 | (OP==`EOR_abx & T==`Ttwo & phi2)
			 | (OP==`EOR_abx & T==`Tthree & phi1)
			 | (OP==`EOR_abx & T==`Tthree & phi2)
			 | (OP==`EOR_abx & T==`Tfour & phi1)
			 | (OP==`LSR_abx & T==`Tzero & phi2)
			 | (OP==`LSR_abx & T==`Tone & phi1)
			 | (OP==`LSR_abx & T==`Ttwo & phi2)
			 | (OP==`LSR_abx & T==`Tthree & phi1)
			 | (OP==`LSR_abx & T==`Tthree & phi2)
			 | (OP==`LSR_abx & T==`Tfour & phi1)
			 | (OP==`LSR_abx & T==`Tfive & phi2)
			 | (OP==`LSR_abx & T==`Tsix & phi1)
			 | (OP==`RTS & T==`Tzero & phi1)
			 | (OP==`RTS & T==`Tzero & phi2)
			 | (OP==`RTS & T==`Tone & phi1)
			 | (OP==`RTS & T==`Tone & phi2)
			 | (OP==`RTS & T==`Ttwo & phi2)
			 | (OP==`RTS & T==`Tthree & phi1)
			 | (OP==`RTS & T==`Tthree & phi2)
			 | (OP==`RTS & T==`Tfour & phi1)
			 | (OP==`RTS & T==`Tfour & phi2)
			 | (OP==`RTS & T==`Tfive & phi1)
			 | (OP==`RTS & T==`Tfive & phi2)
			 | (OP==`ADC_izx & T==`Tzero & phi2)
			 | (OP==`ADC_izx & T==`Tone & phi1)
			 | (OP==`ADC_izx & T==`Tthree & phi2)
			 | (OP==`ADC_izx & T==`Tfour & phi1)
			 | (OP==`ADC_izx & T==`Tfour & phi2)
			 | (OP==`ADC_izx & T==`Tfive & phi1)
			 | (OP==`ADC_zp & T==`Tzero & phi2)
			 | (OP==`ADC_zp & T==`Tone & phi1)
			 | (OP==`ROR_zp & T==`Tzero & phi2)
			 | (OP==`ROR_zp & T==`Tone & phi1)
			 | (OP==`ROR_zp & T==`Tthree & phi2)
			 | (OP==`ROR_zp & T==`Tfour & phi1)
			 | (OP==`PLA & T==`Tzero & phi1)
			 | (OP==`PLA & T==`Tzero & phi2)
			 | (OP==`PLA & T==`Tone & phi1)
			 | (OP==`PLA & T==`Tone & phi2)
			 | (OP==`PLA & T==`Ttwo & phi2)
			 | (OP==`PLA & T==`Tthree & phi1)
			 | (OP==`PLA & T==`Tthree & phi2)
			 | (OP==`ADC_imm & T==`Tone & phi1)
			 | (OP==`ADC_imm & T==`Ttwo & phi2)
			 | (OP==`JMP_zp & T==`Tzero & phi1)
			 | (OP==`JMP_zp & T==`Tzero & phi2)
			 | (OP==`JMP_zp & T==`Tone & phi1)
			 | (OP==`JMP_zp & T==`Ttwo & phi2)
			 | (OP==`JMP_zp & T==`Tthree & phi1)
			 | (OP==`JMP_zp & T==`Tfour & phi2)
			 | (OP==`ADC_abs & T==`Tzero & phi2)
			 | (OP==`ADC_abs & T==`Tone & phi1)
			 | (OP==`ADC_abs & T==`Ttwo & phi2)
			 | (OP==`ADC_abs & T==`Tthree & phi1)
			 | (OP==`ROR_abs & T==`Tzero & phi2)
			 | (OP==`ROR_abs & T==`Tone & phi1)
			 | (OP==`ROR_abs & T==`Ttwo & phi2)
			 | (OP==`ROR_abs & T==`Tthree & phi1)
			 | (OP==`ROR_abs & T==`Tfour & phi2)
			 | (OP==`ROR_abs & T==`Tfive & phi1)
			 | (OP==`BVS_rel & T==`Tzero & phi2)
			 | (OP==`BVS_rel & T==`Ttwo & phi2)
			 | (OP==`BVS_rel & T==`Tthree & phi1)
			 | (OP==`BVS_rel & T==`T1BranchCross & phi1)
			 | (OP==`BVS_rel & T==`T1NoBranch & phi1)
			 | (OP==`ADC_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ADC_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`ADC_izy & T==`TzeroCrossPg & phi2)
			 | (OP==`ADC_izy & T==`Tone & phi1)
			 | (OP==`ADC_izy & T==`Ttwo & phi2)
			 | (OP==`ADC_izy & T==`Tthree & phi1)
			 | (OP==`ADC_izy & T==`Tthree & phi2)
			 | (OP==`ADC_izy & T==`Tfour & phi1)
			 | (OP==`ADC_izy & T==`Tfour & phi2)
			 | (OP==`ADC_izy & T==`Tfive & phi1)
			 | (OP==`ADC_zpx & T==`Tzero & phi2)
			 | (OP==`ADC_zpx & T==`Tone & phi1)
			 | (OP==`ROR_zpx & T==`Tzero & phi2)
			 | (OP==`ROR_zpx & T==`Tone & phi1)
			 | (OP==`ROR_zpx & T==`Tfour & phi2)
			 | (OP==`ROR_zpx & T==`Tfive & phi1)
			 | (OP==`ADC_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ADC_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`ADC_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`ADC_aby & T==`Tone & phi1)
			 | (OP==`ADC_aby & T==`Ttwo & phi2)
			 | (OP==`ADC_aby & T==`Tthree & phi1)
			 | (OP==`ADC_aby & T==`Tthree & phi2)
			 | (OP==`ADC_aby & T==`Tfour & phi1)
			 | (OP==`ADC_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ADC_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`ADC_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`ADC_abx & T==`Tone & phi1)
			 | (OP==`ADC_abx & T==`Ttwo & phi2)
			 | (OP==`ADC_abx & T==`Tthree & phi1)
			 | (OP==`ADC_abx & T==`Tthree & phi2)
			 | (OP==`ADC_abx & T==`Tfour & phi1)
			 | (OP==`ROR_abx & T==`Tzero & phi2)
			 | (OP==`ROR_abx & T==`Tone & phi1)
			 | (OP==`ROR_abx & T==`Ttwo & phi2)
			 | (OP==`ROR_abx & T==`Tthree & phi1)
			 | (OP==`ROR_abx & T==`Tthree & phi2)
			 | (OP==`ROR_abx & T==`Tfour & phi1)
			 | (OP==`ROR_abx & T==`Tfive & phi2)
			 | (OP==`ROR_abx & T==`Tsix & phi1)
			 | (OP==`STA_izx & T==`Tzero & phi2)
			 | (OP==`STA_izx & T==`Tone & phi1)
			 | (OP==`STA_izx & T==`Tthree & phi2)
			 | (OP==`STA_izx & T==`Tfour & phi1)
			 | (OP==`STA_izx & T==`Tfour & phi2)
			 | (OP==`STA_izx & T==`Tfive & phi1)
			 | (OP==`STY_zp & T==`Tzero & phi2)
			 | (OP==`STY_zp & T==`Tone & phi1)
			 | (OP==`STA_zp & T==`Tzero & phi2)
			 | (OP==`STA_zp & T==`Tone & phi1)
			 | (OP==`STX_zp & T==`Tzero & phi2)
			 | (OP==`STX_zp & T==`Tone & phi1)
			 | (OP==`STY_abs & T==`Tzero & phi2)
			 | (OP==`STY_abs & T==`Tone & phi1)
			 | (OP==`STY_abs & T==`Ttwo & phi2)
			 | (OP==`STY_abs & T==`Tthree & phi1)
			 | (OP==`STA_abs & T==`Tzero & phi2)
			 | (OP==`STA_abs & T==`Tone & phi1)
			 | (OP==`STA_abs & T==`Ttwo & phi2)
			 | (OP==`STA_abs & T==`Tthree & phi1)
			 | (OP==`STX_abs & T==`Tzero & phi2)
			 | (OP==`STX_abs & T==`Tone & phi1)
			 | (OP==`STX_abs & T==`Ttwo & phi2)
			 | (OP==`STX_abs & T==`Tthree & phi1)
			 | (OP==`BCC_rel & T==`Tzero & phi2)
			 | (OP==`BCC_rel & T==`Ttwo & phi2)
			 | (OP==`BCC_rel & T==`Tthree & phi1)
			 | (OP==`BCC_rel & T==`T1BranchCross & phi1)
			 | (OP==`BCC_rel & T==`T1NoBranch & phi1)
			 | (OP==`STA_izy & T==`Tzero & phi2)
			 | (OP==`STA_izy & T==`Tone & phi1)
			 | (OP==`STA_izy & T==`Ttwo & phi2)
			 | (OP==`STA_izy & T==`Tthree & phi1)
			 | (OP==`STA_izy & T==`Tthree & phi2)
			 | (OP==`STA_izy & T==`Tfour & phi1)
			 | (OP==`STA_izy & T==`Tfour & phi2)
			 | (OP==`STA_izy & T==`Tfive & phi1)
			 | (OP==`STY_zpx & T==`Tzero & phi2)
			 | (OP==`STY_zpx & T==`Tone & phi1)
			 | (OP==`STA_zpx & T==`Tzero & phi2)
			 | (OP==`STA_zpx & T==`Tone & phi1)
			 | (OP==`STX_zpy & T==`Tzero & phi2)
			 | (OP==`STX_zpy & T==`Tone & phi1)
			 | (OP==`STA_aby & T==`Tzero & phi2)
			 | (OP==`STA_aby & T==`Tone & phi1)
			 | (OP==`STA_aby & T==`Ttwo & phi2)
			 | (OP==`STA_aby & T==`Tthree & phi1)
			 | (OP==`STA_aby & T==`Tthree & phi2)
			 | (OP==`STA_aby & T==`Tfour & phi1)
			 | (OP==`STA_abx & T==`Tzero & phi2)
			 | (OP==`STA_abx & T==`Tone & phi1)
			 | (OP==`STA_abx & T==`Ttwo & phi2)
			 | (OP==`STA_abx & T==`Tthree & phi1)
			 | (OP==`STA_abx & T==`Tthree & phi2)
			 | (OP==`STA_abx & T==`Tfour & phi1)
			 | (OP==`LDY_imm & T==`Tone & phi1)
			 | (OP==`LDY_imm & T==`Ttwo & phi2)
			 | (OP==`LDA_izx & T==`Tzero & phi2)
			 | (OP==`LDA_izx & T==`Tone & phi1)
			 | (OP==`LDA_izx & T==`Tthree & phi2)
			 | (OP==`LDA_izx & T==`Tfour & phi1)
			 | (OP==`LDA_izx & T==`Tfour & phi2)
			 | (OP==`LDA_izx & T==`Tfive & phi1)
			 | (OP==`LDX_imm & T==`Tone & phi1)
			 | (OP==`LDX_imm & T==`Ttwo & phi2)
			 | (OP==`LDY_zp & T==`Tzero & phi2)
			 | (OP==`LDY_zp & T==`Tone & phi1)
			 | (OP==`LDA_zp & T==`Tzero & phi2)
			 | (OP==`LDA_zp & T==`Tone & phi1)
			 | (OP==`LDX_zp & T==`Tzero & phi2)
			 | (OP==`LDX_zp & T==`Tone & phi1)
			 | (OP==`LDA_imm & T==`Tone & phi1)
			 | (OP==`LDA_imm & T==`Ttwo & phi2)
			 | (OP==`LDY_abs & T==`Tzero & phi2)
			 | (OP==`LDY_abs & T==`Tone & phi1)
			 | (OP==`LDY_abs & T==`Ttwo & phi2)
			 | (OP==`LDY_abs & T==`Tthree & phi1)
			 | (OP==`LDA_abs & T==`Tzero & phi2)
			 | (OP==`LDA_abs & T==`Tone & phi1)
			 | (OP==`LDA_abs & T==`Ttwo & phi2)
			 | (OP==`LDA_abs & T==`Tthree & phi1)
			 | (OP==`LDX_abs & T==`Tzero & phi2)
			 | (OP==`LDX_abs & T==`Tone & phi1)
			 | (OP==`LDX_abs & T==`Ttwo & phi2)
			 | (OP==`LDX_abs & T==`Tthree & phi1)
			 | (OP==`BCS_rel & T==`Tzero & phi2)
			 | (OP==`BCS_rel & T==`Ttwo & phi2)
			 | (OP==`BCS_rel & T==`Tthree & phi1)
			 | (OP==`BCS_rel & T==`T1BranchCross & phi1)
			 | (OP==`BCS_rel & T==`T1NoBranch & phi1)
			 | (OP==`LDA_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDA_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`LDA_izy & T==`TzeroCrossPg & phi2)
			 | (OP==`LDA_izy & T==`Tone & phi1)
			 | (OP==`LDA_izy & T==`Ttwo & phi2)
			 | (OP==`LDA_izy & T==`Tthree & phi1)
			 | (OP==`LDA_izy & T==`Tthree & phi2)
			 | (OP==`LDA_izy & T==`Tfour & phi1)
			 | (OP==`LDA_izy & T==`Tfour & phi2)
			 | (OP==`LDA_izy & T==`Tfive & phi1)
			 | (OP==`LDY_zpx & T==`Tzero & phi2)
			 | (OP==`LDY_zpx & T==`Tone & phi1)
			 | (OP==`LDA_zpx & T==`Tzero & phi2)
			 | (OP==`LDA_zpx & T==`Tone & phi1)
			 | (OP==`LDX_zpy & T==`Tzero & phi2)
			 | (OP==`LDX_zpy & T==`Tone & phi1)
			 | (OP==`LDA_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDA_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`LDA_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`LDA_aby & T==`Tone & phi1)
			 | (OP==`LDA_aby & T==`Ttwo & phi2)
			 | (OP==`LDA_aby & T==`Tthree & phi1)
			 | (OP==`LDA_aby & T==`Tthree & phi2)
			 | (OP==`LDA_aby & T==`Tfour & phi1)
			 | (OP==`LDY_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDY_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`LDY_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`LDY_abx & T==`Tone & phi1)
			 | (OP==`LDY_abx & T==`Ttwo & phi2)
			 | (OP==`LDY_abx & T==`Tthree & phi1)
			 | (OP==`LDY_abx & T==`Tthree & phi2)
			 | (OP==`LDY_abx & T==`Tfour & phi1)
			 | (OP==`LDA_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDA_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`LDA_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`LDA_abx & T==`Tone & phi1)
			 | (OP==`LDA_abx & T==`Ttwo & phi2)
			 | (OP==`LDA_abx & T==`Tthree & phi1)
			 | (OP==`LDA_abx & T==`Tthree & phi2)
			 | (OP==`LDA_abx & T==`Tfour & phi1)
			 | (OP==`LDX_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDX_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`LDX_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`LDX_aby & T==`Tone & phi1)
			 | (OP==`LDX_aby & T==`Ttwo & phi2)
			 | (OP==`LDX_aby & T==`Tthree & phi1)
			 | (OP==`LDX_aby & T==`Tthree & phi2)
			 | (OP==`LDX_aby & T==`Tfour & phi1)
			 | (OP==`CPY_imm & T==`Tone & phi1)
			 | (OP==`CPY_imm & T==`Ttwo & phi2)
			 | (OP==`CMP_izx & T==`Tzero & phi2)
			 | (OP==`CMP_izx & T==`Tone & phi1)
			 | (OP==`CMP_izx & T==`Tthree & phi2)
			 | (OP==`CMP_izx & T==`Tfour & phi1)
			 | (OP==`CMP_izx & T==`Tfour & phi2)
			 | (OP==`CMP_izx & T==`Tfive & phi1)
			 | (OP==`CPY_zp & T==`Tzero & phi2)
			 | (OP==`CPY_zp & T==`Tone & phi1)
			 | (OP==`CMP_zp & T==`Tzero & phi2)
			 | (OP==`CMP_zp & T==`Tone & phi1)
			 | (OP==`DEC_zp & T==`Tzero & phi2)
			 | (OP==`DEC_zp & T==`Tone & phi1)
			 | (OP==`DEC_zp & T==`Tthree & phi2)
			 | (OP==`DEC_zp & T==`Tfour & phi1)
			 | (OP==`CMP_imm & T==`Tone & phi1)
			 | (OP==`CMP_imm & T==`Ttwo & phi2)
			 | (OP==`CPY_abs & T==`Tzero & phi2)
			 | (OP==`CPY_abs & T==`Tone & phi1)
			 | (OP==`CPY_abs & T==`Ttwo & phi2)
			 | (OP==`CPY_abs & T==`Tthree & phi1)
			 | (OP==`CMP_abs & T==`Tzero & phi2)
			 | (OP==`CMP_abs & T==`Tone & phi1)
			 | (OP==`CMP_abs & T==`Ttwo & phi2)
			 | (OP==`CMP_abs & T==`Tthree & phi1)
			 | (OP==`DEC_abs & T==`Tzero & phi2)
			 | (OP==`DEC_abs & T==`Tone & phi1)
			 | (OP==`DEC_abs & T==`Ttwo & phi2)
			 | (OP==`DEC_abs & T==`Tthree & phi1)
			 | (OP==`DEC_abs & T==`Tfour & phi2)
			 | (OP==`DEC_abs & T==`Tfive & phi1)
			 | (OP==`BNE_rel & T==`Tzero & phi2)
			 | (OP==`BNE_rel & T==`Ttwo & phi2)
			 | (OP==`BNE_rel & T==`Tthree & phi1)
			 | (OP==`BNE_rel & T==`T1BranchCross & phi1)
			 | (OP==`BNE_rel & T==`T1NoBranch & phi1)
			 | (OP==`CMP_izy & T==`TzeroCrossPg & phi2)
			 | (OP==`CMP_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`CMP_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`CMP_izy & T==`Tone & phi1)
			 | (OP==`CMP_izy & T==`Ttwo & phi2)
			 | (OP==`CMP_izy & T==`Tthree & phi1)
			 | (OP==`CMP_izy & T==`Tthree & phi2)
			 | (OP==`CMP_izy & T==`Tfour & phi1)
			 | (OP==`CMP_izy & T==`Tfour & phi2)
			 | (OP==`CMP_izy & T==`Tfive & phi1)
			 | (OP==`CMP_zpx & T==`Tzero & phi2)
			 | (OP==`CMP_zpx & T==`Tone & phi1)
			 | (OP==`DEC_zpx & T==`Tzero & phi2)
			 | (OP==`DEC_zpx & T==`Tone & phi1)
			 | (OP==`DEC_zpx & T==`Tfour & phi2)
			 | (OP==`DEC_zpx & T==`Tfive & phi1)
			 | (OP==`CMP_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`CMP_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`CMP_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`CMP_aby & T==`Tone & phi1)
			 | (OP==`CMP_aby & T==`Ttwo & phi2)
			 | (OP==`CMP_aby & T==`Tthree & phi1)
			 | (OP==`CMP_aby & T==`Tthree & phi2)
			 | (OP==`CMP_aby & T==`Tfour & phi1)
			 | (OP==`CMP_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`CMP_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`CMP_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`CMP_abx & T==`Tone & phi1)
			 | (OP==`CMP_abx & T==`Ttwo & phi2)
			 | (OP==`CMP_abx & T==`Tthree & phi1)
			 | (OP==`CMP_abx & T==`Tthree & phi2)
			 | (OP==`CMP_abx & T==`Tfour & phi1)
			 | (OP==`DEC_abx & T==`Tzero & phi2)
			 | (OP==`DEC_abx & T==`Tone & phi1)
			 | (OP==`DEC_abx & T==`Ttwo & phi2)
			 | (OP==`DEC_abx & T==`Tthree & phi1)
			 | (OP==`DEC_abx & T==`Tthree & phi2)
			 | (OP==`DEC_abx & T==`Tfour & phi1)
			 | (OP==`DEC_abx & T==`Tfive & phi2)
			 | (OP==`DEC_abx & T==`Tsix & phi1)
			 | (OP==`CPX_imm & T==`Tone & phi1)
			 | (OP==`CPX_imm & T==`Ttwo & phi2)
			 | (OP==`SBC_izx & T==`Tzero & phi2)
			 | (OP==`SBC_izx & T==`Tone & phi1)
			 | (OP==`SBC_izx & T==`Tthree & phi2)
			 | (OP==`SBC_izx & T==`Tfour & phi1)
			 | (OP==`SBC_izx & T==`Tfour & phi2)
			 | (OP==`SBC_izx & T==`Tfive & phi1)
			 | (OP==`CPX_zp & T==`Tzero & phi2)
			 | (OP==`CPX_zp & T==`Tone & phi1)
			 | (OP==`SBC_zp & T==`Tzero & phi2)
			 | (OP==`SBC_zp & T==`Tone & phi1)
			 | (OP==`INC_zp & T==`Tzero & phi2)
			 | (OP==`INC_zp & T==`Tone & phi1)
			 | (OP==`INC_zp & T==`Tthree & phi2)
			 | (OP==`INC_zp & T==`Tfour & phi1)
			 | (OP==`SBC_imm & T==`Tone & phi1)
			 | (OP==`SBC_imm & T==`Ttwo & phi2)
			 | (OP==`CPX_abs & T==`Tzero & phi2)
			 | (OP==`CPX_abs & T==`Tone & phi1)
			 | (OP==`CPX_abs & T==`Ttwo & phi2)
			 | (OP==`CPX_abs & T==`Tthree & phi1)
			 | (OP==`SBC_abs & T==`Tzero & phi2)
			 | (OP==`SBC_abs & T==`Tone & phi1)
			 | (OP==`SBC_abs & T==`Ttwo & phi2)
			 | (OP==`SBC_abs & T==`Tthree & phi1)
			 | (OP==`INC_abs & T==`Tzero & phi2)
			 | (OP==`INC_abs & T==`Tone & phi1)
			 | (OP==`INC_abs & T==`Ttwo & phi2)
			 | (OP==`INC_abs & T==`Tthree & phi1)
			 | (OP==`INC_abs & T==`Tfour & phi2)
			 | (OP==`INC_abs & T==`Tfive & phi1)
			 | (OP==`BEQ_rel & T==`Tzero & phi2)
			 | (OP==`BEQ_rel & T==`Ttwo & phi2)
			 | (OP==`BEQ_rel & T==`Tthree & phi1)
			 | (OP==`BEQ_rel & T==`T1BranchCross & phi1)
			 | (OP==`BEQ_rel & T==`T1NoBranch & phi1)
			 | (OP==`SBC_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`SBC_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`SBC_izy & T==`TzeroCrossPg & phi2)
			 | (OP==`SBC_izy & T==`Tone & phi1)
			 | (OP==`SBC_izy & T==`Ttwo & phi2)
			 | (OP==`SBC_izy & T==`Tthree & phi1)
			 | (OP==`SBC_izy & T==`Tthree & phi2)
			 | (OP==`SBC_izy & T==`Tfour & phi1)
			 | (OP==`SBC_izy & T==`Tfour & phi2)
			 | (OP==`SBC_izy & T==`Tfive & phi1)
			 | (OP==`SBC_zpx & T==`Tzero & phi2)
			 | (OP==`SBC_zpx & T==`Tone & phi1)
			 | (OP==`INC_zpx & T==`Tzero & phi2)
			 | (OP==`INC_zpx & T==`Tone & phi1)
			 | (OP==`INC_zpx & T==`Tfour & phi2)
			 | (OP==`INC_zpx & T==`Tfive & phi1)
			 | (OP==`SBC_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`SBC_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`SBC_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`SBC_aby & T==`Tone & phi1)
			 | (OP==`SBC_aby & T==`Ttwo & phi2)
			 | (OP==`SBC_aby & T==`Tthree & phi1)
			 | (OP==`SBC_aby & T==`Tthree & phi2)
			 | (OP==`SBC_aby & T==`Tfour & phi1)
			 | (OP==`SBC_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`SBC_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`SBC_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`SBC_abx & T==`Tone & phi1)
			 | (OP==`SBC_abx & T==`Ttwo & phi2)
			 | (OP==`SBC_abx & T==`Tthree & phi1)
			 | (OP==`SBC_abx & T==`Tthree & phi2)
			 | (OP==`SBC_abx & T==`Tfour & phi1)
			 | (OP==`INC_abx & T==`Tzero & phi2)
			 | (OP==`INC_abx & T==`Tone & phi1)
			 | (OP==`INC_abx & T==`Ttwo & phi2)
			 | (OP==`INC_abx & T==`Tthree & phi1)
			 | (OP==`INC_abx & T==`Tthree & phi2)
			 | (OP==`INC_abx & T==`Tfour & phi1)
			 | (OP==`INC_abx & T==`Tfive & phi2)
			 | (OP==`INC_abx & T==`Tsix & phi1)
			;

assign control[`DL_ADL] = (OP==`ORA_izx & T==`Ttwo & phi2)
			 | (OP==`ORA_izx & T==`Tthree & phi1)
			 | (OP==`ORA_zp & T==`Tzero & phi1)
			 | (OP==`ORA_zp & T==`Ttwo & phi2)
			 | (OP==`ASL_zp & T==`Ttwo & phi2)
			 | (OP==`ASL_zp & T==`Tthree & phi1)
			 | (OP==`ORA_izy & T==`Ttwo & phi2)
			 | (OP==`ORA_izy & T==`Tthree & phi1)
			 | (OP==`ORA_zpx & T==`Ttwo & phi2)
			 | (OP==`ORA_zpx & T==`Tthree & phi1)
			 | (OP==`ASL_zpx & T==`Ttwo & phi2)
			 | (OP==`ASL_zpx & T==`Tthree & phi1)
			 | (OP==`AND_izx & T==`Ttwo & phi2)
			 | (OP==`AND_izx & T==`Tthree & phi1)
			 | (OP==`BIT_zp & T==`Tzero & phi1)
			 | (OP==`BIT_zp & T==`Ttwo & phi2)
			 | (OP==`AND_zp & T==`Tzero & phi1)
			 | (OP==`AND_zp & T==`Ttwo & phi2)
			 | (OP==`ROL_zp & T==`Ttwo & phi2)
			 | (OP==`ROL_zp & T==`Tthree & phi1)
			 | (OP==`AND_izy & T==`Ttwo & phi2)
			 | (OP==`AND_izy & T==`Tthree & phi1)
			 | (OP==`AND_zpx & T==`Ttwo & phi2)
			 | (OP==`AND_zpx & T==`Tthree & phi1)
			 | (OP==`ROL_zpx & T==`Ttwo & phi2)
			 | (OP==`ROL_zpx & T==`Tthree & phi1)
			 | (OP==`EOR_izx & T==`Ttwo & phi2)
			 | (OP==`EOR_izx & T==`Tthree & phi1)
			 | (OP==`EOR_zp & T==`Tzero & phi1)
			 | (OP==`EOR_zp & T==`Ttwo & phi2)
			 | (OP==`LSR_zp & T==`Ttwo & phi2)
			 | (OP==`LSR_zp & T==`Tthree & phi1)
			 | (OP==`EOR_izy & T==`Ttwo & phi2)
			 | (OP==`EOR_izy & T==`Tthree & phi1)
			 | (OP==`EOR_zpx & T==`Ttwo & phi2)
			 | (OP==`EOR_zpx & T==`Tthree & phi1)
			 | (OP==`LSR_zpx & T==`Ttwo & phi2)
			 | (OP==`LSR_zpx & T==`Tthree & phi1)
			 | (OP==`ADC_izx & T==`Ttwo & phi2)
			 | (OP==`ADC_izx & T==`Tthree & phi1)
			 | (OP==`ADC_zp & T==`Tzero & phi1)
			 | (OP==`ADC_zp & T==`Ttwo & phi2)
			 | (OP==`ROR_zp & T==`Ttwo & phi2)
			 | (OP==`ROR_zp & T==`Tthree & phi1)
			 | (OP==`ADC_izy & T==`Ttwo & phi2)
			 | (OP==`ADC_izy & T==`Tthree & phi1)
			 | (OP==`ADC_zpx & T==`Ttwo & phi2)
			 | (OP==`ADC_zpx & T==`Tthree & phi1)
			 | (OP==`ROR_zpx & T==`Ttwo & phi2)
			 | (OP==`ROR_zpx & T==`Tthree & phi1)
			 | (OP==`STA_izx & T==`Ttwo & phi2)
			 | (OP==`STA_izx & T==`Tthree & phi1)
			 | (OP==`STY_zp & T==`Tzero & phi1)
			 | (OP==`STY_zp & T==`Ttwo & phi2)
			 | (OP==`STA_zp & T==`Tzero & phi1)
			 | (OP==`STA_zp & T==`Ttwo & phi2)
			 | (OP==`STX_zp & T==`Tzero & phi1)
			 | (OP==`STX_zp & T==`Ttwo & phi2)
			 | (OP==`STA_izy & T==`Ttwo & phi2)
			 | (OP==`STA_izy & T==`Tthree & phi1)
			 | (OP==`STY_zpx & T==`Ttwo & phi2)
			 | (OP==`STY_zpx & T==`Tthree & phi1)
			 | (OP==`STA_zpx & T==`Ttwo & phi2)
			 | (OP==`STA_zpx & T==`Tthree & phi1)
			 | (OP==`STX_zpy & T==`Ttwo & phi2)
			 | (OP==`STX_zpy & T==`Tthree & phi1)
			 | (OP==`LDA_izx & T==`Ttwo & phi2)
			 | (OP==`LDA_izx & T==`Tthree & phi1)
			 | (OP==`LDY_zp & T==`Tzero & phi1)
			 | (OP==`LDY_zp & T==`Ttwo & phi2)
			 | (OP==`LDA_zp & T==`Tzero & phi1)
			 | (OP==`LDA_zp & T==`Ttwo & phi2)
			 | (OP==`LDX_zp & T==`Tzero & phi1)
			 | (OP==`LDX_zp & T==`Ttwo & phi2)
			 | (OP==`LDA_izy & T==`Ttwo & phi2)
			 | (OP==`LDA_izy & T==`Tthree & phi1)
			 | (OP==`LDY_zpx & T==`Ttwo & phi2)
			 | (OP==`LDY_zpx & T==`Tthree & phi1)
			 | (OP==`LDA_zpx & T==`Ttwo & phi2)
			 | (OP==`LDA_zpx & T==`Tthree & phi1)
			 | (OP==`LDX_zpy & T==`Ttwo & phi2)
			 | (OP==`LDX_zpy & T==`Tthree & phi1)
			 | (OP==`CMP_izx & T==`Ttwo & phi2)
			 | (OP==`CMP_izx & T==`Tthree & phi1)
			 | (OP==`CPY_zp & T==`Tzero & phi1)
			 | (OP==`CPY_zp & T==`Ttwo & phi2)
			 | (OP==`CMP_zp & T==`Tzero & phi1)
			 | (OP==`CMP_zp & T==`Ttwo & phi2)
			 | (OP==`DEC_zp & T==`Ttwo & phi2)
			 | (OP==`DEC_zp & T==`Tthree & phi1)
			 | (OP==`CMP_izy & T==`Ttwo & phi2)
			 | (OP==`CMP_izy & T==`Tthree & phi1)
			 | (OP==`CMP_zpx & T==`Ttwo & phi2)
			 | (OP==`CMP_zpx & T==`Tthree & phi1)
			 | (OP==`DEC_zpx & T==`Ttwo & phi2)
			 | (OP==`DEC_zpx & T==`Tthree & phi1)
			 | (OP==`SBC_izx & T==`Ttwo & phi2)
			 | (OP==`SBC_izx & T==`Tthree & phi1)
			 | (OP==`CPX_zp & T==`Tzero & phi1)
			 | (OP==`CPX_zp & T==`Ttwo & phi2)
			 | (OP==`SBC_zp & T==`Tzero & phi1)
			 | (OP==`SBC_zp & T==`Ttwo & phi2)
			 | (OP==`INC_zp & T==`Ttwo & phi2)
			 | (OP==`INC_zp & T==`Tthree & phi1)
			 | (OP==`SBC_izy & T==`Ttwo & phi2)
			 | (OP==`SBC_izy & T==`Tthree & phi1)
			 | (OP==`SBC_zpx & T==`Ttwo & phi2)
			 | (OP==`SBC_zpx & T==`Tthree & phi1)
			 | (OP==`INC_zpx & T==`Ttwo & phi2)
			 | (OP==`INC_zpx & T==`Tthree & phi1)
			;

assign control[`DL_ADH] = (OP==`BRK & T==`Tzero & phi2)
			 | (OP==`BRK & T==`Tone & phi1)
			 | (OP==`ORA_izx & T==`Tzero & phi1)
			 | (OP==`ORA_izx & T==`Tfive & phi2)
			 | (OP==`ORA_abs & T==`Tzero & phi1)
			 | (OP==`ORA_abs & T==`Tthree & phi2)
			 | (OP==`ASL_abs & T==`Tthree & phi2)
			 | (OP==`ASL_abs & T==`Tfour & phi1)
			 | (OP==`ORA_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ORA_izy & T==`Tfour & phi2)
			 | (OP==`ORA_izy & T==`Tfive & phi1)
			 | (OP==`ORA_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ORA_aby & T==`Tthree & phi2)
			 | (OP==`ORA_aby & T==`Tfour & phi1)
			 | (OP==`ORA_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ORA_abx & T==`Tthree & phi2)
			 | (OP==`ORA_abx & T==`Tfour & phi1)
			 | (OP==`ASL_abx & T==`Tthree & phi2)
			 | (OP==`ASL_abx & T==`Tfour & phi1)
			 | (OP==`JSR_abs & T==`Tzero & phi2)
			 | (OP==`JSR_abs & T==`Tone & phi1)
			 | (OP==`AND_izx & T==`Tzero & phi1)
			 | (OP==`AND_izx & T==`Tfive & phi2)
			 | (OP==`BIT_abs & T==`Tzero & phi1)
			 | (OP==`BIT_abs & T==`Tthree & phi2)
			 | (OP==`AND_abs & T==`Tzero & phi1)
			 | (OP==`AND_abs & T==`Tthree & phi2)
			 | (OP==`ROL_abs & T==`Tthree & phi2)
			 | (OP==`ROL_abs & T==`Tfour & phi1)
			 | (OP==`AND_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`AND_izy & T==`Tfour & phi2)
			 | (OP==`AND_izy & T==`Tfive & phi1)
			 | (OP==`AND_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`AND_aby & T==`Tthree & phi2)
			 | (OP==`AND_aby & T==`Tfour & phi1)
			 | (OP==`AND_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`AND_abx & T==`Tthree & phi2)
			 | (OP==`AND_abx & T==`Tfour & phi1)
			 | (OP==`ROL_abx & T==`Tthree & phi2)
			 | (OP==`ROL_abx & T==`Tfour & phi1)
			 | (OP==`RTI & T==`Tzero & phi2)
			 | (OP==`RTI & T==`Tone & phi1)
			 | (OP==`EOR_izx & T==`Tzero & phi1)
			 | (OP==`EOR_izx & T==`Tfive & phi2)
			 | (OP==`JMP_abs & T==`Tzero & phi2)
			 | (OP==`JMP_abs & T==`Tone & phi1)
			 | (OP==`EOR_abs & T==`Tzero & phi1)
			 | (OP==`EOR_abs & T==`Tthree & phi2)
			 | (OP==`LSR_abs & T==`Tthree & phi2)
			 | (OP==`LSR_abs & T==`Tfour & phi1)
			 | (OP==`EOR_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`EOR_izy & T==`Tfour & phi2)
			 | (OP==`EOR_izy & T==`Tfive & phi1)
			 | (OP==`EOR_aby & T==`Tthree & phi2)
			 | (OP==`EOR_aby & T==`Tfour & phi1)
			 | (OP==`EOR_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`EOR_abx & T==`Tthree & phi2)
			 | (OP==`EOR_abx & T==`Tfour & phi1)
			 | (OP==`LSR_abx & T==`Tthree & phi2)
			 | (OP==`LSR_abx & T==`Tfour & phi1)
			 | (OP==`RTS & T==`Tzero & phi1)
			 | (OP==`RTS & T==`Tfive & phi2)
			 | (OP==`ADC_izx & T==`Tzero & phi1)
			 | (OP==`ADC_izx & T==`Tfive & phi2)
			 | (OP==`JMP_zp & T==`Tzero & phi2)
			 | (OP==`JMP_zp & T==`Tone & phi1)
			 | (OP==`JMP_zp & T==`Tthree & phi2)
			 | (OP==`JMP_zp & T==`Tfour & phi1)
			 | (OP==`ADC_abs & T==`Tzero & phi1)
			 | (OP==`ADC_abs & T==`Tthree & phi2)
			 | (OP==`ROR_abs & T==`Tthree & phi2)
			 | (OP==`ROR_abs & T==`Tfour & phi1)
			 | (OP==`ADC_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ADC_izy & T==`Tfour & phi2)
			 | (OP==`ADC_izy & T==`Tfive & phi1)
			 | (OP==`ADC_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ADC_aby & T==`Tthree & phi2)
			 | (OP==`ADC_aby & T==`Tfour & phi1)
			 | (OP==`ADC_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ADC_abx & T==`Tthree & phi2)
			 | (OP==`ADC_abx & T==`Tfour & phi1)
			 | (OP==`ROR_abx & T==`Tthree & phi2)
			 | (OP==`ROR_abx & T==`Tfour & phi1)
			 | (OP==`STA_izx & T==`Tzero & phi1)
			 | (OP==`STA_izx & T==`Tfive & phi2)
			 | (OP==`STY_abs & T==`Tzero & phi1)
			 | (OP==`STY_abs & T==`Tthree & phi2)
			 | (OP==`STA_abs & T==`Tzero & phi1)
			 | (OP==`STA_abs & T==`Tthree & phi2)
			 | (OP==`STX_abs & T==`Tzero & phi1)
			 | (OP==`STX_abs & T==`Tthree & phi2)
			 | (OP==`STA_izy & T==`Tfour & phi2)
			 | (OP==`STA_izy & T==`Tfive & phi1)
			 | (OP==`STA_aby & T==`Tthree & phi2)
			 | (OP==`STA_aby & T==`Tfour & phi1)
			 | (OP==`STA_abx & T==`Tthree & phi2)
			 | (OP==`STA_abx & T==`Tfour & phi1)
			 | (OP==`LDA_izx & T==`Tzero & phi1)
			 | (OP==`LDA_izx & T==`Tfive & phi2)
			 | (OP==`LDY_abs & T==`Tzero & phi1)
			 | (OP==`LDY_abs & T==`Tthree & phi2)
			 | (OP==`LDA_abs & T==`Tzero & phi1)
			 | (OP==`LDA_abs & T==`Tthree & phi2)
			 | (OP==`LDX_abs & T==`Tzero & phi1)
			 | (OP==`LDX_abs & T==`Tthree & phi2)
			 | (OP==`LDA_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDA_izy & T==`Tfour & phi2)
			 | (OP==`LDA_izy & T==`Tfive & phi1)
			 | (OP==`LDA_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDA_aby & T==`Tthree & phi2)
			 | (OP==`LDA_aby & T==`Tfour & phi1)
			 | (OP==`LDY_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDY_abx & T==`Tthree & phi2)
			 | (OP==`LDY_abx & T==`Tfour & phi1)
			 | (OP==`LDA_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDA_abx & T==`Tthree & phi2)
			 | (OP==`LDA_abx & T==`Tfour & phi1)
			 | (OP==`LDX_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDX_aby & T==`Tthree & phi2)
			 | (OP==`LDX_aby & T==`Tfour & phi1)
			 | (OP==`CMP_izx & T==`Tzero & phi1)
			 | (OP==`CMP_izx & T==`Tfive & phi2)
			 | (OP==`CPY_abs & T==`Tzero & phi1)
			 | (OP==`CPY_abs & T==`Tthree & phi2)
			 | (OP==`CMP_abs & T==`Tzero & phi1)
			 | (OP==`CMP_abs & T==`Tthree & phi2)
			 | (OP==`DEC_abs & T==`Tthree & phi2)
			 | (OP==`DEC_abs & T==`Tfour & phi1)
			 | (OP==`CMP_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`CMP_izy & T==`Tfour & phi2)
			 | (OP==`CMP_izy & T==`Tfive & phi1)
			 | (OP==`CMP_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`CMP_aby & T==`Tthree & phi2)
			 | (OP==`CMP_aby & T==`Tfour & phi1)
			 | (OP==`CMP_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`CMP_abx & T==`Tthree & phi2)
			 | (OP==`CMP_abx & T==`Tfour & phi1)
			 | (OP==`DEC_abx & T==`Tthree & phi2)
			 | (OP==`DEC_abx & T==`Tfour & phi1)
			 | (OP==`SBC_izx & T==`Tzero & phi1)
			 | (OP==`SBC_izx & T==`Tfive & phi2)
			 | (OP==`CPX_abs & T==`Tzero & phi1)
			 | (OP==`CPX_abs & T==`Tthree & phi2)
			 | (OP==`SBC_abs & T==`Tzero & phi1)
			 | (OP==`SBC_abs & T==`Tthree & phi2)
			 | (OP==`INC_abs & T==`Tthree & phi2)
			 | (OP==`INC_abs & T==`Tfour & phi1)
			 | (OP==`SBC_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`SBC_izy & T==`Tfour & phi2)
			 | (OP==`SBC_izy & T==`Tfive & phi1)
			 | (OP==`SBC_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`SBC_aby & T==`Tthree & phi2)
			 | (OP==`SBC_aby & T==`Tfour & phi1)
			 | (OP==`SBC_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`SBC_abx & T==`Tthree & phi2)
			 | (OP==`SBC_abx & T==`Tfour & phi1)
			 | (OP==`INC_abx & T==`Tthree & phi2)
			 | (OP==`INC_abx & T==`Tfour & phi1)
			;

assign control[`O_ADH0] = (OP==`ORA_izx & T==`Ttwo & phi2)
			 | (OP==`ORA_izx & T==`Tthree & phi1)
			 | (OP==`ORA_zp & T==`Tzero & phi1)
			 | (OP==`ORA_zp & T==`Ttwo & phi2)
			 | (OP==`ASL_zp & T==`Ttwo & phi2)
			 | (OP==`ASL_zp & T==`Tthree & phi1)
			 | (OP==`ORA_izy & T==`Ttwo & phi2)
			 | (OP==`ORA_izy & T==`Tthree & phi1)
			 | (OP==`ORA_zpx & T==`Ttwo & phi2)
			 | (OP==`ORA_zpx & T==`Tthree & phi1)
			 | (OP==`ASL_zpx & T==`Ttwo & phi2)
			 | (OP==`ASL_zpx & T==`Tthree & phi1)
			 | (OP==`AND_izx & T==`Ttwo & phi2)
			 | (OP==`AND_izx & T==`Tthree & phi1)
			 | (OP==`BIT_zp & T==`Tzero & phi1)
			 | (OP==`BIT_zp & T==`Ttwo & phi2)
			 | (OP==`AND_zp & T==`Tzero & phi1)
			 | (OP==`AND_zp & T==`Ttwo & phi2)
			 | (OP==`ROL_zp & T==`Ttwo & phi2)
			 | (OP==`ROL_zp & T==`Tthree & phi1)
			 | (OP==`AND_izy & T==`Ttwo & phi2)
			 | (OP==`AND_izy & T==`Tthree & phi1)
			 | (OP==`AND_zpx & T==`Ttwo & phi2)
			 | (OP==`AND_zpx & T==`Tthree & phi1)
			 | (OP==`ROL_zpx & T==`Ttwo & phi2)
			 | (OP==`ROL_zpx & T==`Tthree & phi1)
			 | (OP==`EOR_izx & T==`Ttwo & phi2)
			 | (OP==`EOR_izx & T==`Tthree & phi1)
			 | (OP==`EOR_zp & T==`Tzero & phi1)
			 | (OP==`EOR_zp & T==`Ttwo & phi2)
			 | (OP==`LSR_zp & T==`Ttwo & phi2)
			 | (OP==`LSR_zp & T==`Tthree & phi1)
			 | (OP==`EOR_izy & T==`Ttwo & phi2)
			 | (OP==`EOR_izy & T==`Tthree & phi1)
			 | (OP==`EOR_zpx & T==`Ttwo & phi2)
			 | (OP==`EOR_zpx & T==`Tthree & phi1)
			 | (OP==`LSR_zpx & T==`Ttwo & phi2)
			 | (OP==`LSR_zpx & T==`Tthree & phi1)
			 | (OP==`ADC_izx & T==`Ttwo & phi2)
			 | (OP==`ADC_izx & T==`Tthree & phi1)
			 | (OP==`ADC_zp & T==`Tzero & phi1)
			 | (OP==`ADC_zp & T==`Ttwo & phi2)
			 | (OP==`ROR_zp & T==`Ttwo & phi2)
			 | (OP==`ROR_zp & T==`Tthree & phi1)
			 | (OP==`ADC_izy & T==`Ttwo & phi2)
			 | (OP==`ADC_izy & T==`Tthree & phi1)
			 | (OP==`ADC_zpx & T==`Ttwo & phi2)
			 | (OP==`ADC_zpx & T==`Tthree & phi1)
			 | (OP==`ROR_zpx & T==`Ttwo & phi2)
			 | (OP==`ROR_zpx & T==`Tthree & phi1)
			 | (OP==`STA_izx & T==`Ttwo & phi2)
			 | (OP==`STA_izx & T==`Tthree & phi1)
			 | (OP==`STY_zp & T==`Tzero & phi1)
			 | (OP==`STY_zp & T==`Ttwo & phi2)
			 | (OP==`STA_zp & T==`Tzero & phi1)
			 | (OP==`STA_zp & T==`Ttwo & phi2)
			 | (OP==`STX_zp & T==`Tzero & phi1)
			 | (OP==`STX_zp & T==`Ttwo & phi2)
			 | (OP==`STA_izy & T==`Ttwo & phi2)
			 | (OP==`STA_izy & T==`Tthree & phi1)
			 | (OP==`STY_zpx & T==`Ttwo & phi2)
			 | (OP==`STY_zpx & T==`Tthree & phi1)
			 | (OP==`STA_zpx & T==`Ttwo & phi2)
			 | (OP==`STA_zpx & T==`Tthree & phi1)
			 | (OP==`STX_zpy & T==`Ttwo & phi2)
			 | (OP==`STX_zpy & T==`Tthree & phi1)
			 | (OP==`LDA_izx & T==`Ttwo & phi2)
			 | (OP==`LDA_izx & T==`Tthree & phi1)
			 | (OP==`LDY_zp & T==`Tzero & phi1)
			 | (OP==`LDY_zp & T==`Ttwo & phi2)
			 | (OP==`LDA_zp & T==`Tzero & phi1)
			 | (OP==`LDA_zp & T==`Ttwo & phi2)
			 | (OP==`LDX_zp & T==`Tzero & phi1)
			 | (OP==`LDX_zp & T==`Ttwo & phi2)
			 | (OP==`LDA_izy & T==`Ttwo & phi2)
			 | (OP==`LDA_izy & T==`Tthree & phi1)
			 | (OP==`LDY_zpx & T==`Ttwo & phi2)
			 | (OP==`LDY_zpx & T==`Tthree & phi1)
			 | (OP==`LDA_zpx & T==`Ttwo & phi2)
			 | (OP==`LDA_zpx & T==`Tthree & phi1)
			 | (OP==`LDX_zpy & T==`Ttwo & phi2)
			 | (OP==`LDX_zpy & T==`Tthree & phi1)
			 | (OP==`CMP_izx & T==`Ttwo & phi2)
			 | (OP==`CMP_izx & T==`Tthree & phi1)
			 | (OP==`CPY_zp & T==`Tzero & phi1)
			 | (OP==`CPY_zp & T==`Ttwo & phi2)
			 | (OP==`CMP_zp & T==`Tzero & phi1)
			 | (OP==`CMP_zp & T==`Ttwo & phi2)
			 | (OP==`DEC_zp & T==`Ttwo & phi2)
			 | (OP==`DEC_zp & T==`Tthree & phi1)
			 | (OP==`CMP_izy & T==`Ttwo & phi2)
			 | (OP==`CMP_izy & T==`Tthree & phi1)
			 | (OP==`CMP_zpx & T==`Ttwo & phi2)
			 | (OP==`CMP_zpx & T==`Tthree & phi1)
			 | (OP==`DEC_zpx & T==`Ttwo & phi2)
			 | (OP==`DEC_zpx & T==`Tthree & phi1)
			 | (OP==`SBC_izx & T==`Ttwo & phi2)
			 | (OP==`SBC_izx & T==`Tthree & phi1)
			 | (OP==`CPX_zp & T==`Tzero & phi1)
			 | (OP==`CPX_zp & T==`Ttwo & phi2)
			 | (OP==`SBC_zp & T==`Tzero & phi1)
			 | (OP==`SBC_zp & T==`Ttwo & phi2)
			 | (OP==`INC_zp & T==`Ttwo & phi2)
			 | (OP==`INC_zp & T==`Tthree & phi1)
			 | (OP==`SBC_izy & T==`Ttwo & phi2)
			 | (OP==`SBC_izy & T==`Tthree & phi1)
			 | (OP==`SBC_zpx & T==`Ttwo & phi2)
			 | (OP==`SBC_zpx & T==`Tthree & phi1)
			 | (OP==`INC_zpx & T==`Ttwo & phi2)
			 | (OP==`INC_zpx & T==`Tthree & phi1)
			;

assign control[`O_ADH1to7] = (OP==`BRK & T==`Ttwo & phi2)
			 | (OP==`BRK & T==`Tthree & phi1)
			 | (OP==`ORA_izx & T==`Ttwo & phi2)
			 | (OP==`ORA_izx & T==`Tthree & phi1)
			 | (OP==`ORA_zp & T==`Tzero & phi1)
			 | (OP==`ORA_zp & T==`Ttwo & phi2)
			 | (OP==`ASL_zp & T==`Ttwo & phi2)
			 | (OP==`ASL_zp & T==`Tthree & phi1)
			 | (OP==`PHP & T==`Tzero & phi1)
			 | (OP==`PHP & T==`Ttwo & phi2)
			 | (OP==`ORA_izy & T==`Ttwo & phi2)
			 | (OP==`ORA_izy & T==`Tthree & phi1)
			 | (OP==`ORA_zpx & T==`Ttwo & phi2)
			 | (OP==`ORA_zpx & T==`Tthree & phi1)
			 | (OP==`ASL_zpx & T==`Ttwo & phi2)
			 | (OP==`ASL_zpx & T==`Tthree & phi1)
			 | (OP==`JSR_abs & T==`Ttwo & phi2)
			 | (OP==`JSR_abs & T==`Tthree & phi1)
			 | (OP==`AND_izx & T==`Ttwo & phi2)
			 | (OP==`AND_izx & T==`Tthree & phi1)
			 | (OP==`BIT_zp & T==`Tzero & phi1)
			 | (OP==`BIT_zp & T==`Ttwo & phi2)
			 | (OP==`AND_zp & T==`Tzero & phi1)
			 | (OP==`AND_zp & T==`Ttwo & phi2)
			 | (OP==`ROL_zp & T==`Ttwo & phi2)
			 | (OP==`ROL_zp & T==`Tthree & phi1)
			 | (OP==`PLP & T==`Ttwo & phi2)
			 | (OP==`PLP & T==`Tthree & phi1)
			 | (OP==`AND_izy & T==`Ttwo & phi2)
			 | (OP==`AND_izy & T==`Tthree & phi1)
			 | (OP==`AND_zpx & T==`Ttwo & phi2)
			 | (OP==`AND_zpx & T==`Tthree & phi1)
			 | (OP==`ROL_zpx & T==`Ttwo & phi2)
			 | (OP==`ROL_zpx & T==`Tthree & phi1)
			 | (OP==`RTI & T==`Ttwo & phi2)
			 | (OP==`RTI & T==`Tthree & phi1)
			 | (OP==`EOR_izx & T==`Ttwo & phi2)
			 | (OP==`EOR_izx & T==`Tthree & phi1)
			 | (OP==`EOR_zp & T==`Tzero & phi1)
			 | (OP==`EOR_zp & T==`Ttwo & phi2)
			 | (OP==`LSR_zp & T==`Ttwo & phi2)
			 | (OP==`LSR_zp & T==`Tthree & phi1)
			 | (OP==`PHA & T==`Tzero & phi1)
			 | (OP==`PHA & T==`Ttwo & phi2)
			 | (OP==`EOR_izy & T==`Ttwo & phi2)
			 | (OP==`EOR_izy & T==`Tthree & phi1)
			 | (OP==`EOR_zpx & T==`Ttwo & phi2)
			 | (OP==`EOR_zpx & T==`Tthree & phi1)
			 | (OP==`LSR_zpx & T==`Ttwo & phi2)
			 | (OP==`LSR_zpx & T==`Tthree & phi1)
			 | (OP==`RTS & T==`Ttwo & phi2)
			 | (OP==`RTS & T==`Tthree & phi1)
			 | (OP==`ADC_izx & T==`Ttwo & phi2)
			 | (OP==`ADC_izx & T==`Tthree & phi1)
			 | (OP==`ADC_zp & T==`Tzero & phi1)
			 | (OP==`ADC_zp & T==`Ttwo & phi2)
			 | (OP==`ROR_zp & T==`Ttwo & phi2)
			 | (OP==`ROR_zp & T==`Tthree & phi1)
			 | (OP==`PLA & T==`Ttwo & phi2)
			 | (OP==`PLA & T==`Tthree & phi1)
			 | (OP==`ADC_izy & T==`Ttwo & phi2)
			 | (OP==`ADC_izy & T==`Tthree & phi1)
			 | (OP==`ADC_zpx & T==`Ttwo & phi2)
			 | (OP==`ADC_zpx & T==`Tthree & phi1)
			 | (OP==`ROR_zpx & T==`Ttwo & phi2)
			 | (OP==`ROR_zpx & T==`Tthree & phi1)
			 | (OP==`STA_izx & T==`Ttwo & phi2)
			 | (OP==`STA_izx & T==`Tthree & phi1)
			 | (OP==`STY_zp & T==`Tzero & phi1)
			 | (OP==`STY_zp & T==`Ttwo & phi2)
			 | (OP==`STA_zp & T==`Tzero & phi1)
			 | (OP==`STA_zp & T==`Ttwo & phi2)
			 | (OP==`STX_zp & T==`Tzero & phi1)
			 | (OP==`STX_zp & T==`Ttwo & phi2)
			 | (OP==`STA_izy & T==`Ttwo & phi2)
			 | (OP==`STA_izy & T==`Tthree & phi1)
			 | (OP==`STY_zpx & T==`Ttwo & phi2)
			 | (OP==`STY_zpx & T==`Tthree & phi1)
			 | (OP==`STA_zpx & T==`Ttwo & phi2)
			 | (OP==`STA_zpx & T==`Tthree & phi1)
			 | (OP==`STX_zpy & T==`Ttwo & phi2)
			 | (OP==`STX_zpy & T==`Tthree & phi1)
			 | (OP==`LDA_izx & T==`Ttwo & phi2)
			 | (OP==`LDA_izx & T==`Tthree & phi1)
			 | (OP==`LDY_zp & T==`Tzero & phi1)
			 | (OP==`LDY_zp & T==`Ttwo & phi2)
			 | (OP==`LDA_zp & T==`Tzero & phi1)
			 | (OP==`LDA_zp & T==`Ttwo & phi2)
			 | (OP==`LDX_zp & T==`Tzero & phi1)
			 | (OP==`LDX_zp & T==`Ttwo & phi2)
			 | (OP==`LDA_izy & T==`Ttwo & phi2)
			 | (OP==`LDA_izy & T==`Tthree & phi1)
			 | (OP==`LDY_zpx & T==`Ttwo & phi2)
			 | (OP==`LDY_zpx & T==`Tthree & phi1)
			 | (OP==`LDA_zpx & T==`Ttwo & phi2)
			 | (OP==`LDA_zpx & T==`Tthree & phi1)
			 | (OP==`LDX_zpy & T==`Ttwo & phi2)
			 | (OP==`LDX_zpy & T==`Tthree & phi1)
			 | (OP==`CMP_izx & T==`Ttwo & phi2)
			 | (OP==`CMP_izx & T==`Tthree & phi1)
			 | (OP==`CPY_zp & T==`Tzero & phi1)
			 | (OP==`CPY_zp & T==`Ttwo & phi2)
			 | (OP==`CMP_zp & T==`Tzero & phi1)
			 | (OP==`CMP_zp & T==`Ttwo & phi2)
			 | (OP==`DEC_zp & T==`Ttwo & phi2)
			 | (OP==`DEC_zp & T==`Tthree & phi1)
			 | (OP==`CMP_izy & T==`Ttwo & phi2)
			 | (OP==`CMP_izy & T==`Tthree & phi1)
			 | (OP==`CMP_zpx & T==`Ttwo & phi2)
			 | (OP==`CMP_zpx & T==`Tthree & phi1)
			 | (OP==`DEC_zpx & T==`Ttwo & phi2)
			 | (OP==`DEC_zpx & T==`Tthree & phi1)
			 | (OP==`SBC_izx & T==`Ttwo & phi2)
			 | (OP==`SBC_izx & T==`Tthree & phi1)
			 | (OP==`CPX_zp & T==`Tzero & phi1)
			 | (OP==`CPX_zp & T==`Ttwo & phi2)
			 | (OP==`SBC_zp & T==`Tzero & phi1)
			 | (OP==`SBC_zp & T==`Ttwo & phi2)
			 | (OP==`INC_zp & T==`Ttwo & phi2)
			 | (OP==`INC_zp & T==`Tthree & phi1)
			 | (OP==`SBC_izy & T==`Ttwo & phi2)
			 | (OP==`SBC_izy & T==`Tthree & phi1)
			 | (OP==`SBC_zpx & T==`Ttwo & phi2)
			 | (OP==`SBC_zpx & T==`Tthree & phi1)
			 | (OP==`INC_zpx & T==`Ttwo & phi2)
			 | (OP==`INC_zpx & T==`Tthree & phi1)
			;

assign control[`nADH_ABH] = (OP==`BRK & T==`Tzero & phi1)
			 | (OP==`BRK & T==`Tthree & phi2)
			 | (OP==`BRK & T==`Tfour & phi1)
			 | (OP==`BRK & T==`Tfour & phi2)
			 | (OP==`BRK & T==`Tfive & phi1)
			 | (OP==`BRK & T==`Tsix & phi2)
			 | (OP==`ORA_izx & T==`Tthree & phi2)
			 | (OP==`ORA_izx & T==`Tfour & phi1)
			 | (OP==`ORA_izx & T==`Tfour & phi2)
			 | (OP==`ORA_izx & T==`Tfive & phi1)
			 | (OP==`ASL_zp & T==`Tzero & phi1)
			 | (OP==`ASL_zp & T==`Tthree & phi2)
			 | (OP==`ASL_zp & T==`Tfour & phi1)
			 | (OP==`ASL_zp & T==`Tfour & phi2)
			 | (OP==`ASL_abs & T==`Tzero & phi1)
			 | (OP==`ASL_abs & T==`Tfour & phi2)
			 | (OP==`ASL_abs & T==`Tfive & phi1)
			 | (OP==`ASL_abs & T==`Tfive & phi2)
			 | (OP==`BPL_rel & T==`Tzero & phi1)
			 | (OP==`BPL_rel & T==`Tthree & phi2)
			 | (OP==`BPL_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`ORA_izy & T==`Tthree & phi2)
			 | (OP==`ORA_izy & T==`Tfour & phi1)
			 | (OP==`ORA_zpx & T==`Tzero & phi1)
			 | (OP==`ORA_zpx & T==`Tthree & phi2)
			 | (OP==`ASL_zpx & T==`Tzero & phi1)
			 | (OP==`ASL_zpx & T==`Tthree & phi2)
			 | (OP==`ASL_zpx & T==`Tfour & phi1)
			 | (OP==`ASL_zpx & T==`Tfour & phi2)
			 | (OP==`ASL_zpx & T==`Tfive & phi1)
			 | (OP==`ASL_zpx & T==`Tfive & phi2)
			 | (OP==`ASL_abx & T==`Tzero & phi1)
			 | (OP==`ASL_abx & T==`Tfour & phi2 & !carry)
			 | (OP==`ASL_abx & T==`Tfive & phi1)
			 | (OP==`ASL_abx & T==`Tfive & phi2)
			 | (OP==`ASL_abx & T==`Tsix & phi1)
			 | (OP==`ASL_abx & T==`Tsix & phi2)
			 | (OP==`JSR_abs & T==`Tthree & phi2)
			 | (OP==`JSR_abs & T==`Tfour & phi1)
			 | (OP==`JSR_abs & T==`Tfour & phi2)
			 | (OP==`JSR_abs & T==`Tfive & phi1)
			 | (OP==`AND_izx & T==`Tthree & phi2)
			 | (OP==`AND_izx & T==`Tfour & phi1)
			 | (OP==`AND_izx & T==`Tfour & phi2)
			 | (OP==`AND_izx & T==`Tfive & phi1)
			 | (OP==`ROL_zp & T==`Tzero & phi1)
			 | (OP==`ROL_zp & T==`Tthree & phi2)
			 | (OP==`ROL_zp & T==`Tfour & phi1)
			 | (OP==`ROL_zp & T==`Tfour & phi2)
			 | (OP==`PLP & T==`Tzero & phi1)
			 | (OP==`PLP & T==`Tthree & phi2)
			 | (OP==`ROL_abs & T==`Tzero & phi1)
			 | (OP==`ROL_abs & T==`Tfour & phi2)
			 | (OP==`ROL_abs & T==`Tfive & phi1)
			 | (OP==`ROL_abs & T==`Tfive & phi2)
			 | (OP==`BMI_rel & T==`Tzero & phi1)
			 | (OP==`BMI_rel & T==`Tthree & phi2)
			 | (OP==`BMI_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`AND_izy & T==`Tthree & phi2)
			 | (OP==`AND_izy & T==`Tfour & phi1)
			 | (OP==`AND_zpx & T==`Tzero & phi1)
			 | (OP==`AND_zpx & T==`Tthree & phi2)
			 | (OP==`ROL_zpx & T==`Tzero & phi1)
			 | (OP==`ROL_zpx & T==`Tthree & phi2)
			 | (OP==`ROL_zpx & T==`Tfour & phi1)
			 | (OP==`ROL_zpx & T==`Tfour & phi2)
			 | (OP==`ROL_zpx & T==`Tfive & phi1)
			 | (OP==`ROL_zpx & T==`Tfive & phi2)
			 | (OP==`ROL_abx & T==`Tzero & phi1)
			 | (OP==`ROL_abx & T==`Tfour & phi2 & !carry)
			 | (OP==`ROL_abx & T==`Tfive & phi1)
			 | (OP==`ROL_abx & T==`Tfive & phi2)
			 | (OP==`ROL_abx & T==`Tsix & phi1)
			 | (OP==`ROL_abx & T==`Tsix & phi2)
			 | (OP==`RTI & T==`Tzero & phi1)
			 | (OP==`RTI & T==`Tthree & phi2)
			 | (OP==`RTI & T==`Tfour & phi1)
			 | (OP==`RTI & T==`Tfour & phi2)
			 | (OP==`RTI & T==`Tfive & phi1)
			 | (OP==`RTI & T==`Tfive & phi2)
			 | (OP==`EOR_izx & T==`Tthree & phi2)
			 | (OP==`EOR_izx & T==`Tfour & phi1)
			 | (OP==`EOR_izx & T==`Tfour & phi2)
			 | (OP==`EOR_izx & T==`Tfive & phi1)
			 | (OP==`LSR_zp & T==`Tzero & phi1)
			 | (OP==`LSR_zp & T==`Tthree & phi2)
			 | (OP==`LSR_zp & T==`Tfour & phi1)
			 | (OP==`LSR_zp & T==`Tfour & phi2)
			 | (OP==`LSR_abs & T==`Tzero & phi1)
			 | (OP==`LSR_abs & T==`Tfour & phi2)
			 | (OP==`LSR_abs & T==`Tfive & phi1)
			 | (OP==`LSR_abs & T==`Tfive & phi2)
			 | (OP==`BVC_rel & T==`Tzero & phi1)
			 | (OP==`BVC_rel & T==`Tthree & phi2)
			 | (OP==`BVC_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`EOR_izy & T==`Tthree & phi2)
			 | (OP==`EOR_izy & T==`Tfour & phi1)
			 | (OP==`EOR_zpx & T==`Tzero & phi1)
			 | (OP==`EOR_zpx & T==`Tthree & phi2)
			 | (OP==`LSR_zpx & T==`Tzero & phi1)
			 | (OP==`LSR_zpx & T==`Tthree & phi2)
			 | (OP==`LSR_zpx & T==`Tfour & phi1)
			 | (OP==`LSR_zpx & T==`Tfour & phi2)
			 | (OP==`LSR_zpx & T==`Tfive & phi1)
			 | (OP==`LSR_zpx & T==`Tfive & phi2)
			 | (OP==`LSR_abx & T==`Tzero & phi1)
			 | (OP==`LSR_abx & T==`Tfour & phi2 & !carry)
			 | (OP==`LSR_abx & T==`Tfive & phi1)
			 | (OP==`LSR_abx & T==`Tfive & phi2)
			 | (OP==`LSR_abx & T==`Tsix & phi1)
			 | (OP==`LSR_abx & T==`Tsix & phi2)
			 | (OP==`RTS & T==`Tthree & phi2)
			 | (OP==`RTS & T==`Tfour & phi1)
			 | (OP==`RTS & T==`Tfour & phi2)
			 | (OP==`RTS & T==`Tfive & phi1)
			 | (OP==`ADC_izx & T==`Tthree & phi2)
			 | (OP==`ADC_izx & T==`Tfour & phi1)
			 | (OP==`ADC_izx & T==`Tfour & phi2)
			 | (OP==`ADC_izx & T==`Tfive & phi1)
			 | (OP==`ROR_zp & T==`Tzero & phi1)
			 | (OP==`ROR_zp & T==`Tthree & phi2)
			 | (OP==`ROR_zp & T==`Tfour & phi1)
			 | (OP==`ROR_zp & T==`Tfour & phi2)
			 | (OP==`PLA & T==`Tzero & phi1)
			 | (OP==`PLA & T==`Tthree & phi2)
			 | (OP==`JMP_zp & T==`Tzero & phi1)
			 | (OP==`JMP_zp & T==`Tfour & phi2)
			 | (OP==`ROR_abs & T==`Tzero & phi1)
			 | (OP==`ROR_abs & T==`Tfour & phi2)
			 | (OP==`ROR_abs & T==`Tfive & phi1)
			 | (OP==`ROR_abs & T==`Tfive & phi2)
			 | (OP==`BVS_rel & T==`Tzero & phi1)
			 | (OP==`BVS_rel & T==`Tthree & phi2)
			 | (OP==`BVS_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`ADC_izy & T==`Tthree & phi2)
			 | (OP==`ADC_izy & T==`Tfour & phi1)
			 | (OP==`ADC_zpx & T==`Tzero & phi1)
			 | (OP==`ADC_zpx & T==`Tthree & phi2)
			 | (OP==`ROR_zpx & T==`Tzero & phi1)
			 | (OP==`ROR_zpx & T==`Tthree & phi2)
			 | (OP==`ROR_zpx & T==`Tfour & phi1)
			 | (OP==`ROR_zpx & T==`Tfour & phi2)
			 | (OP==`ROR_zpx & T==`Tfive & phi1)
			 | (OP==`ROR_zpx & T==`Tfive & phi2)
			 | (OP==`ROR_abx & T==`Tzero & phi1)
			 | (OP==`ROR_abx & T==`Tfour & phi2 & !carry)
			 | (OP==`ROR_abx & T==`Tfive & phi1)
			 | (OP==`ROR_abx & T==`Tfive & phi2)
			 | (OP==`ROR_abx & T==`Tsix & phi1)
			 | (OP==`ROR_abx & T==`Tsix & phi2)
			 | (OP==`STA_izx & T==`Tthree & phi2)
			 | (OP==`STA_izx & T==`Tfour & phi1)
			 | (OP==`STA_izx & T==`Tfour & phi2)
			 | (OP==`STA_izx & T==`Tfive & phi1)
			 | (OP==`BCC_rel & T==`Tzero & phi1)
			 | (OP==`BCC_rel & T==`Tthree & phi2)
			 | (OP==`BCC_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`STA_izy & T==`Tzero & phi1)
			 | (OP==`STA_izy & T==`Tthree & phi2)
			 | (OP==`STA_izy & T==`Tfour & phi1)
			 | (OP==`STA_izy & T==`Tfive & phi2 & !carry)
			 | (OP==`STY_zpx & T==`Tzero & phi1)
			 | (OP==`STY_zpx & T==`Tthree & phi2)
			 | (OP==`STA_zpx & T==`Tzero & phi1)
			 | (OP==`STA_zpx & T==`Tthree & phi2)
			 | (OP==`STX_zpy & T==`Tzero & phi1)
			 | (OP==`STX_zpy & T==`Tthree & phi2)
			 | (OP==`STA_aby & T==`Tzero & phi1)
			 | (OP==`STA_aby & T==`Tfour & phi2 & !carry)
			 | (OP==`STA_abx & T==`Tzero & phi1)
			 | (OP==`STA_abx & T==`Tfour & phi2 & !carry)
			 | (OP==`LDA_izx & T==`Tthree & phi2)
			 | (OP==`LDA_izx & T==`Tfour & phi1)
			 | (OP==`LDA_izx & T==`Tfour & phi2)
			 | (OP==`LDA_izx & T==`Tfive & phi1)
			 | (OP==`BCS_rel & T==`Tzero & phi1)
			 | (OP==`BCS_rel & T==`Tthree & phi2)
			 | (OP==`BCS_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`LDA_izy & T==`Tthree & phi2)
			 | (OP==`LDA_izy & T==`Tfour & phi1)
			 | (OP==`LDY_zpx & T==`Tzero & phi1)
			 | (OP==`LDY_zpx & T==`Tthree & phi2)
			 | (OP==`LDA_zpx & T==`Tzero & phi1)
			 | (OP==`LDA_zpx & T==`Tthree & phi2)
			 | (OP==`LDX_zpy & T==`Tzero & phi1)
			 | (OP==`LDX_zpy & T==`Tthree & phi2)
			 | (OP==`CMP_izx & T==`Tthree & phi2)
			 | (OP==`CMP_izx & T==`Tfour & phi1)
			 | (OP==`CMP_izx & T==`Tfour & phi2)
			 | (OP==`CMP_izx & T==`Tfive & phi1)
			 | (OP==`DEC_zp & T==`Tzero & phi1)
			 | (OP==`DEC_zp & T==`Tthree & phi2)
			 | (OP==`DEC_zp & T==`Tfour & phi1)
			 | (OP==`DEC_zp & T==`Tfour & phi2)
			 | (OP==`DEC_abs & T==`Tzero & phi1)
			 | (OP==`DEC_abs & T==`Tfour & phi2)
			 | (OP==`DEC_abs & T==`Tfive & phi1)
			 | (OP==`DEC_abs & T==`Tfive & phi2)
			 | (OP==`BNE_rel & T==`Tzero & phi1)
			 | (OP==`BNE_rel & T==`Tthree & phi2)
			 | (OP==`BNE_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`CMP_izy & T==`Tthree & phi2)
			 | (OP==`CMP_izy & T==`Tfour & phi1)
			 | (OP==`CMP_zpx & T==`Tzero & phi1)
			 | (OP==`CMP_zpx & T==`Tthree & phi2)
			 | (OP==`DEC_zpx & T==`Tzero & phi1)
			 | (OP==`DEC_zpx & T==`Tthree & phi2)
			 | (OP==`DEC_zpx & T==`Tfour & phi1)
			 | (OP==`DEC_zpx & T==`Tfour & phi2)
			 | (OP==`DEC_zpx & T==`Tfive & phi1)
			 | (OP==`DEC_zpx & T==`Tfive & phi2)
			 | (OP==`DEC_abx & T==`Tzero & phi1)
			 | (OP==`DEC_abx & T==`Tfour & phi2 & !carry)
			 | (OP==`DEC_abx & T==`Tfive & phi1)
			 | (OP==`DEC_abx & T==`Tfive & phi2)
			 | (OP==`DEC_abx & T==`Tsix & phi1)
			 | (OP==`DEC_abx & T==`Tsix & phi2)
			 | (OP==`SBC_izx & T==`Tthree & phi2)
			 | (OP==`SBC_izx & T==`Tfour & phi1)
			 | (OP==`SBC_izx & T==`Tfour & phi2)
			 | (OP==`SBC_izx & T==`Tfive & phi1)
			 | (OP==`INC_zp & T==`Tzero & phi1)
			 | (OP==`INC_zp & T==`Tthree & phi2)
			 | (OP==`INC_zp & T==`Tfour & phi1)
			 | (OP==`INC_zp & T==`Tfour & phi2)
			 | (OP==`INC_abs & T==`Tzero & phi1)
			 | (OP==`INC_abs & T==`Tfour & phi2)
			 | (OP==`INC_abs & T==`Tfive & phi1)
			 | (OP==`INC_abs & T==`Tfive & phi2)
			 | (OP==`BEQ_rel & T==`Tzero & phi1)
			 | (OP==`BEQ_rel & T==`Tthree & phi2)
			 | (OP==`BEQ_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`SBC_izy & T==`Tthree & phi2)
			 | (OP==`SBC_izy & T==`Tfour & phi1)
			 | (OP==`SBC_zpx & T==`Tzero & phi1)
			 | (OP==`SBC_zpx & T==`Tthree & phi2)
			 | (OP==`INC_zpx & T==`Tzero & phi1)
			 | (OP==`INC_zpx & T==`Tthree & phi2)
			 | (OP==`INC_zpx & T==`Tfour & phi1)
			 | (OP==`INC_zpx & T==`Tfour & phi2)
			 | (OP==`INC_zpx & T==`Tfive & phi1)
			 | (OP==`INC_zpx & T==`Tfive & phi2)
			 | (OP==`INC_abx & T==`Tzero & phi1)
			 | (OP==`INC_abx & T==`Tfour & phi2 & !carry)
			 | (OP==`INC_abx & T==`Tfive & phi1)
			 | (OP==`INC_abx & T==`Tfive & phi2)
			 | (OP==`INC_abx & T==`Tsix & phi1)
			 | (OP==`INC_abx & T==`Tsix & phi2)
			;

assign control[`nADL_ABL] = (OP==`ASL_zp & T==`Tzero & phi1)
			 | (OP==`ASL_zp & T==`Tthree & phi2)
			 | (OP==`ASL_zp & T==`Tfour & phi1)
			 | (OP==`ASL_zp & T==`Tfour & phi2)
			 | (OP==`ASL_abs & T==`Tzero & phi1)
			 | (OP==`ASL_abs & T==`Tfour & phi2)
			 | (OP==`ASL_abs & T==`Tfive & phi1)
			 | (OP==`ASL_abs & T==`Tfive & phi2)
			 | (OP==`ORA_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`ORA_izy & T==`Tfive & phi2)
			 | (OP==`ASL_zpx & T==`Tzero & phi1)
			 | (OP==`ASL_zpx & T==`Tfour & phi2)
			 | (OP==`ASL_zpx & T==`Tfive & phi1)
			 | (OP==`ASL_zpx & T==`Tfive & phi2)
			 | (OP==`ORA_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`ORA_aby & T==`Tfour & phi2)
			 | (OP==`ORA_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`ORA_abx & T==`Tfour & phi2)
			 | (OP==`ASL_abx & T==`Tzero & phi1)
			 | (OP==`ASL_abx & T==`Tfour & phi2)
			 | (OP==`ASL_abx & T==`Tfive & phi1)
			 | (OP==`ASL_abx & T==`Tfive & phi2)
			 | (OP==`ASL_abx & T==`Tsix & phi1)
			 | (OP==`ASL_abx & T==`Tsix & phi2)
			 | (OP==`ROL_zp & T==`Tzero & phi1)
			 | (OP==`ROL_zp & T==`Tthree & phi2)
			 | (OP==`ROL_zp & T==`Tfour & phi1)
			 | (OP==`ROL_zp & T==`Tfour & phi2)
			 | (OP==`ROL_abs & T==`Tzero & phi1)
			 | (OP==`ROL_abs & T==`Tfour & phi2)
			 | (OP==`ROL_abs & T==`Tfive & phi1)
			 | (OP==`ROL_abs & T==`Tfive & phi2)
			 | (OP==`AND_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`AND_izy & T==`Tfive & phi2)
			 | (OP==`ROL_zpx & T==`Tzero & phi1)
			 | (OP==`ROL_zpx & T==`Tfour & phi2)
			 | (OP==`ROL_zpx & T==`Tfive & phi1)
			 | (OP==`ROL_zpx & T==`Tfive & phi2)
			 | (OP==`AND_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`AND_aby & T==`Tfour & phi2)
			 | (OP==`AND_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`AND_abx & T==`Tfour & phi2)
			 | (OP==`ROL_abx & T==`Tzero & phi1)
			 | (OP==`ROL_abx & T==`Tfour & phi2)
			 | (OP==`ROL_abx & T==`Tfive & phi1)
			 | (OP==`ROL_abx & T==`Tfive & phi2)
			 | (OP==`ROL_abx & T==`Tsix & phi1)
			 | (OP==`ROL_abx & T==`Tsix & phi2)
			 | (OP==`LSR_zp & T==`Tzero & phi1)
			 | (OP==`LSR_zp & T==`Tthree & phi2)
			 | (OP==`LSR_zp & T==`Tfour & phi1)
			 | (OP==`LSR_zp & T==`Tfour & phi2)
			 | (OP==`LSR_abs & T==`Tzero & phi1)
			 | (OP==`LSR_abs & T==`Tfour & phi2)
			 | (OP==`LSR_abs & T==`Tfive & phi1)
			 | (OP==`LSR_abs & T==`Tfive & phi2)
			 | (OP==`EOR_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`EOR_izy & T==`Tfive & phi2)
			 | (OP==`LSR_zpx & T==`Tzero & phi1)
			 | (OP==`LSR_zpx & T==`Tfour & phi2)
			 | (OP==`LSR_zpx & T==`Tfive & phi1)
			 | (OP==`LSR_zpx & T==`Tfive & phi2)
			 | (OP==`EOR_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`EOR_aby & T==`Tfour & phi2)
			 | (OP==`EOR_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`EOR_abx & T==`Tfour & phi2)
			 | (OP==`LSR_abx & T==`Tzero & phi1)
			 | (OP==`LSR_abx & T==`Tfour & phi2)
			 | (OP==`LSR_abx & T==`Tfive & phi1)
			 | (OP==`LSR_abx & T==`Tfive & phi2)
			 | (OP==`LSR_abx & T==`Tsix & phi1)
			 | (OP==`LSR_abx & T==`Tsix & phi2)
			 | (OP==`ROR_zp & T==`Tzero & phi1)
			 | (OP==`ROR_zp & T==`Tthree & phi2)
			 | (OP==`ROR_zp & T==`Tfour & phi1)
			 | (OP==`ROR_zp & T==`Tfour & phi2)
			 | (OP==`ROR_abs & T==`Tzero & phi1)
			 | (OP==`ROR_abs & T==`Tfour & phi2)
			 | (OP==`ROR_abs & T==`Tfive & phi1)
			 | (OP==`ROR_abs & T==`Tfive & phi2)
			 | (OP==`ADC_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`ADC_izy & T==`Tfive & phi2)
			 | (OP==`ROR_zpx & T==`Tzero & phi1)
			 | (OP==`ROR_zpx & T==`Tfour & phi2)
			 | (OP==`ROR_zpx & T==`Tfive & phi1)
			 | (OP==`ROR_zpx & T==`Tfive & phi2)
			 | (OP==`ADC_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`ADC_aby & T==`Tfour & phi1)
			 | (OP==`ADC_aby & T==`Tfour & phi2)
			 | (OP==`ROR_abx & T==`Tzero & phi1)
			 | (OP==`ROR_abx & T==`Tfour & phi2)
			 | (OP==`ROR_abx & T==`Tfive & phi1)
			 | (OP==`ROR_abx & T==`Tfive & phi2)
			 | (OP==`ROR_abx & T==`Tsix & phi1)
			 | (OP==`ROR_abx & T==`Tsix & phi2)
			 | (OP==`STA_izy & T==`Tzero & phi1)
			 | (OP==`STA_izy & T==`Tfive & phi2)
			 | (OP==`STA_aby & T==`Tzero & phi1)
			 | (OP==`STA_aby & T==`Tfour & phi2)
			 | (OP==`STA_abx & T==`Tzero & phi1)
			 | (OP==`STA_abx & T==`Tfour & phi2)
			 | (OP==`LDA_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`LDA_izy & T==`Tfive & phi2)
			 | (OP==`LDA_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`LDA_aby & T==`Tfour & phi2)
			 | (OP==`LDY_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`LDY_abx & T==`Tfour & phi2)
			 | (OP==`LDA_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`LDA_abx & T==`Tfour & phi2)
			 | (OP==`LDX_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`LDX_aby & T==`Tfour & phi2)
			 | (OP==`DEC_zp & T==`Tzero & phi1)
			 | (OP==`DEC_zp & T==`Tthree & phi2)
			 | (OP==`DEC_zp & T==`Tfour & phi1)
			 | (OP==`DEC_zp & T==`Tfour & phi2)
			 | (OP==`DEC_abs & T==`Tzero & phi1)
			 | (OP==`DEC_abs & T==`Tfour & phi2)
			 | (OP==`DEC_abs & T==`Tfive & phi1)
			 | (OP==`DEC_abs & T==`Tfive & phi2)
			 | (OP==`CMP_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`CMP_izy & T==`Tfive & phi2)
			 | (OP==`DEC_zpx & T==`Tzero & phi1)
			 | (OP==`DEC_zpx & T==`Tfour & phi2)
			 | (OP==`DEC_zpx & T==`Tfive & phi1)
			 | (OP==`DEC_zpx & T==`Tfive & phi2)
			 | (OP==`CMP_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`CMP_aby & T==`Tfour & phi2)
			 | (OP==`CMP_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`CMP_abx & T==`Tfour & phi2)
			 | (OP==`DEC_abx & T==`Tzero & phi1)
			 | (OP==`DEC_abx & T==`Tfour & phi2)
			 | (OP==`DEC_abx & T==`Tfive & phi1)
			 | (OP==`DEC_abx & T==`Tfive & phi2)
			 | (OP==`DEC_abx & T==`Tsix & phi1)
			 | (OP==`DEC_abx & T==`Tsix & phi2)
			 | (OP==`INC_zp & T==`Tzero & phi1)
			 | (OP==`INC_zp & T==`Tthree & phi2)
			 | (OP==`INC_zp & T==`Tfour & phi1)
			 | (OP==`INC_zp & T==`Tfour & phi2)
			 | (OP==`INC_abs & T==`Tzero & phi1)
			 | (OP==`INC_abs & T==`Tfour & phi2)
			 | (OP==`INC_abs & T==`Tfive & phi1)
			 | (OP==`INC_abs & T==`Tfive & phi2)
			 | (OP==`SBC_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`SBC_izy & T==`Tfive & phi2)
			 | (OP==`INC_zpx & T==`Tzero & phi1)
			 | (OP==`INC_zpx & T==`Tfour & phi2)
			 | (OP==`INC_zpx & T==`Tfive & phi1)
			 | (OP==`INC_zpx & T==`Tfive & phi2)
			 | (OP==`SBC_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`SBC_aby & T==`Tfour & phi2)
			 | (OP==`SBC_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`SBC_abx & T==`Tfour & phi2)
			 | (OP==`INC_abx & T==`Tzero & phi1)
			 | (OP==`INC_abx & T==`Tfour & phi2)
			 | (OP==`INC_abx & T==`Tfive & phi1)
			 | (OP==`INC_abx & T==`Tfive & phi2)
			 | (OP==`INC_abx & T==`Tsix & phi1)
			 | (OP==`INC_abx & T==`Tsix & phi2)
			;

assign control[`PCL_PCL] = (OP==`BRK & T==`Tzero & phi1)
			 | (OP==`BRK & T==`Tthree & phi1)
			 | (OP==`BRK & T==`Tfour & phi1)
			 | (OP==`BRK & T==`Tfive & phi1)
			 | (OP==`BRK & T==`Tsix & phi1)
			 | (OP==`ORA_izx & T==`Tzero & phi1)
			 | (OP==`ORA_izx & T==`Tthree & phi1)
			 | (OP==`ORA_izx & T==`Tfour & phi1)
			 | (OP==`ORA_izx & T==`Tfive & phi1)
			 | (OP==`ORA_zp & T==`Tzero & phi1)
			 | (OP==`ASL_zp & T==`Tzero & phi1)
			 | (OP==`ASL_zp & T==`Tthree & phi1)
			 | (OP==`ASL_zp & T==`Tfour & phi1)
			 | (OP==`PHP & T==`Tzero & phi1)
			 | (OP==`ORA_abs & T==`Tzero & phi1)
			 | (OP==`ASL_abs & T==`Tzero & phi1)
			 | (OP==`ASL_abs & T==`Tfour & phi1)
			 | (OP==`ASL_abs & T==`Tfive & phi1)
			 | (OP==`ORA_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`ORA_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ORA_izy & T==`Tthree & phi1)
			 | (OP==`ORA_izy & T==`Tfour & phi1)
			 | (OP==`ORA_izy & T==`Tfive & phi1)
			 | (OP==`ORA_zpx & T==`Tzero & phi1)
			 | (OP==`ORA_zpx & T==`Tthree & phi1)
			 | (OP==`ASL_zpx & T==`Tzero & phi1)
			 | (OP==`ASL_zpx & T==`Tthree & phi1)
			 | (OP==`ASL_zpx & T==`Tfour & phi1)
			 | (OP==`ASL_zpx & T==`Tfive & phi1)
			 | (OP==`ORA_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ORA_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`ORA_aby & T==`Tfour & phi1)
			 | (OP==`ORA_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ORA_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`ORA_abx & T==`Tfour & phi1)
			 | (OP==`ASL_abx & T==`Tzero & phi1)
			 | (OP==`ASL_abx & T==`Tfour & phi1)
			 | (OP==`ASL_abx & T==`Tfive & phi1)
			 | (OP==`ASL_abx & T==`Tsix & phi1)
			 | (OP==`JSR_abs & T==`Tthree & phi1)
			 | (OP==`JSR_abs & T==`Tfour & phi1)
			 | (OP==`JSR_abs & T==`Tfive & phi1)
			 | (OP==`AND_izx & T==`Tzero & phi1)
			 | (OP==`AND_izx & T==`Tthree & phi1)
			 | (OP==`AND_izx & T==`Tfour & phi1)
			 | (OP==`AND_izx & T==`Tfive & phi1)
			 | (OP==`BIT_zp & T==`Tzero & phi1)
			 | (OP==`AND_zp & T==`Tzero & phi1)
			 | (OP==`ROL_zp & T==`Tzero & phi1)
			 | (OP==`ROL_zp & T==`Tthree & phi1)
			 | (OP==`ROL_zp & T==`Tfour & phi1)
			 | (OP==`PLP & T==`Tzero & phi1)
			 | (OP==`PLP & T==`Tthree & phi1)
			 | (OP==`BIT_abs & T==`Tzero & phi1)
			 | (OP==`AND_abs & T==`Tzero & phi1)
			 | (OP==`ROL_abs & T==`Tzero & phi1)
			 | (OP==`ROL_abs & T==`Tfour & phi1)
			 | (OP==`ROL_abs & T==`Tfive & phi1)
			 | (OP==`AND_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`AND_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`AND_izy & T==`Tthree & phi1)
			 | (OP==`AND_izy & T==`Tfour & phi1)
			 | (OP==`AND_izy & T==`Tfive & phi1)
			 | (OP==`AND_zpx & T==`Tzero & phi1)
			 | (OP==`AND_zpx & T==`Tthree & phi1)
			 | (OP==`ROL_zpx & T==`Tzero & phi1)
			 | (OP==`ROL_zpx & T==`Tthree & phi1)
			 | (OP==`ROL_zpx & T==`Tfour & phi1)
			 | (OP==`ROL_zpx & T==`Tfive & phi1)
			 | (OP==`AND_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`AND_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`AND_aby & T==`Tfour & phi1)
			 | (OP==`AND_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`AND_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`AND_abx & T==`Tfour & phi1)
			 | (OP==`ROL_abx & T==`Tzero & phi1)
			 | (OP==`ROL_abx & T==`Tfour & phi1)
			 | (OP==`ROL_abx & T==`Tfive & phi1)
			 | (OP==`ROL_abx & T==`Tsix & phi1)
			 | (OP==`RTI & T==`Tzero & phi1)
			 | (OP==`RTI & T==`Tthree & phi1)
			 | (OP==`RTI & T==`Tfour & phi1)
			 | (OP==`RTI & T==`Tfive & phi1)
			 | (OP==`EOR_izx & T==`Tzero & phi1)
			 | (OP==`EOR_izx & T==`Tthree & phi1)
			 | (OP==`EOR_izx & T==`Tfour & phi1)
			 | (OP==`EOR_izx & T==`Tfive & phi1)
			 | (OP==`EOR_zp & T==`Tzero & phi1)
			 | (OP==`LSR_zp & T==`Tzero & phi1)
			 | (OP==`LSR_zp & T==`Tthree & phi1)
			 | (OP==`LSR_zp & T==`Tfour & phi1)
			 | (OP==`PHA & T==`Tzero & phi1)
			 | (OP==`EOR_abs & T==`Tzero & phi1)
			 | (OP==`LSR_abs & T==`Tzero & phi1)
			 | (OP==`LSR_abs & T==`Tfour & phi1)
			 | (OP==`LSR_abs & T==`Tfive & phi1)
			 | (OP==`EOR_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`EOR_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`EOR_izy & T==`Tthree & phi1)
			 | (OP==`EOR_izy & T==`Tfour & phi1)
			 | (OP==`EOR_izy & T==`Tfive & phi1)
			 | (OP==`EOR_zpx & T==`Tzero & phi1)
			 | (OP==`EOR_zpx & T==`Tthree & phi1)
			 | (OP==`LSR_zpx & T==`Tzero & phi1)
			 | (OP==`LSR_zpx & T==`Tthree & phi1)
			 | (OP==`LSR_zpx & T==`Tfour & phi1)
			 | (OP==`LSR_zpx & T==`Tfive & phi1)
			 | (OP==`EOR_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`EOR_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`EOR_aby & T==`Tfour & phi1)
			 | (OP==`EOR_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`EOR_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`EOR_abx & T==`Tfour & phi1)
			 | (OP==`LSR_abx & T==`Tzero & phi1)
			 | (OP==`LSR_abx & T==`Tfour & phi1)
			 | (OP==`LSR_abx & T==`Tfive & phi1)
			 | (OP==`LSR_abx & T==`Tsix & phi1)
			 | (OP==`RTS & T==`Tthree & phi1)
			 | (OP==`RTS & T==`Tfour & phi1)
			 | (OP==`RTS & T==`Tfive & phi1)
			 | (OP==`ADC_izx & T==`Tzero & phi1)
			 | (OP==`ADC_izx & T==`Tthree & phi1)
			 | (OP==`ADC_izx & T==`Tfour & phi1)
			 | (OP==`ADC_izx & T==`Tfive & phi1)
			 | (OP==`ADC_zp & T==`Tzero & phi1)
			 | (OP==`ROR_zp & T==`Tzero & phi1)
			 | (OP==`ROR_zp & T==`Tthree & phi1)
			 | (OP==`ROR_zp & T==`Tfour & phi1)
			 | (OP==`PLA & T==`Tzero & phi1)
			 | (OP==`PLA & T==`Tthree & phi1)
			 | (OP==`JMP_zp & T==`Tzero & phi1)
			 | (OP==`JMP_zp & T==`Tfour & phi1)
			 | (OP==`ADC_abs & T==`Tzero & phi1)
			 | (OP==`ROR_abs & T==`Tzero & phi1)
			 | (OP==`ROR_abs & T==`Tfour & phi1)
			 | (OP==`ROR_abs & T==`Tfive & phi1)
			 | (OP==`ADC_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ADC_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`ADC_izy & T==`Tthree & phi1)
			 | (OP==`ADC_izy & T==`Tfour & phi1)
			 | (OP==`ADC_izy & T==`Tfive & phi1)
			 | (OP==`ADC_zpx & T==`Tzero & phi1)
			 | (OP==`ADC_zpx & T==`Tthree & phi1)
			 | (OP==`ROR_zpx & T==`Tzero & phi1)
			 | (OP==`ROR_zpx & T==`Tthree & phi1)
			 | (OP==`ROR_zpx & T==`Tfour & phi1)
			 | (OP==`ROR_zpx & T==`Tfive & phi1)
			 | (OP==`ADC_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ADC_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`ADC_aby & T==`Tfour & phi1)
			 | (OP==`ADC_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ADC_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`ADC_abx & T==`Tfour & phi1)
			 | (OP==`ROR_abx & T==`Tzero & phi1)
			 | (OP==`ROR_abx & T==`Tfour & phi1)
			 | (OP==`ROR_abx & T==`Tfive & phi1)
			 | (OP==`ROR_abx & T==`Tsix & phi1)
			 | (OP==`STA_izx & T==`Tzero & phi1)
			 | (OP==`STA_izx & T==`Tthree & phi1)
			 | (OP==`STA_izx & T==`Tfour & phi1)
			 | (OP==`STA_izx & T==`Tfive & phi1)
			 | (OP==`STY_zp & T==`Tzero & phi1)
			 | (OP==`STA_zp & T==`Tzero & phi1)
			 | (OP==`STX_zp & T==`Tzero & phi1)
			 | (OP==`STY_abs & T==`Tzero & phi1)
			 | (OP==`STA_abs & T==`Tzero & phi1)
			 | (OP==`STX_abs & T==`Tzero & phi1)
			 | (OP==`STA_izy & T==`Tzero & phi1)
			 | (OP==`STA_izy & T==`Tthree & phi1)
			 | (OP==`STA_izy & T==`Tfour & phi1)
			 | (OP==`STA_izy & T==`Tfive & phi1)
			 | (OP==`STY_zpx & T==`Tzero & phi1)
			 | (OP==`STY_zpx & T==`Tthree & phi1)
			 | (OP==`STA_zpx & T==`Tzero & phi1)
			 | (OP==`STA_zpx & T==`Tthree & phi1)
			 | (OP==`STX_zpy & T==`Tzero & phi1)
			 | (OP==`STX_zpy & T==`Tthree & phi1)
			 | (OP==`STA_aby & T==`Tzero & phi1)
			 | (OP==`STA_aby & T==`Tfour & phi1)
			 | (OP==`STA_abx & T==`Tzero & phi1)
			 | (OP==`STA_abx & T==`Tfour & phi1)
			 | (OP==`LDA_izx & T==`Tzero & phi1)
			 | (OP==`LDA_izx & T==`Tthree & phi1)
			 | (OP==`LDA_izx & T==`Tfour & phi1)
			 | (OP==`LDA_izx & T==`Tfive & phi1)
			 | (OP==`LDY_zp & T==`Tzero & phi1)
			 | (OP==`LDA_zp & T==`Tzero & phi1)
			 | (OP==`LDX_zp & T==`Tzero & phi1)
			 | (OP==`LDY_abs & T==`Tzero & phi1)
			 | (OP==`LDA_abs & T==`Tzero & phi1)
			 | (OP==`LDX_abs & T==`Tzero & phi1)
			 | (OP==`LDA_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDA_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`LDA_izy & T==`Tthree & phi1)
			 | (OP==`LDA_izy & T==`Tfour & phi1)
			 | (OP==`LDA_izy & T==`Tfive & phi1)
			 | (OP==`LDY_zpx & T==`Tzero & phi1)
			 | (OP==`LDY_zpx & T==`Tthree & phi1)
			 | (OP==`LDA_zpx & T==`Tzero & phi1)
			 | (OP==`LDA_zpx & T==`Tthree & phi1)
			 | (OP==`LDX_zpy & T==`Tzero & phi1)
			 | (OP==`LDX_zpy & T==`Tthree & phi1)
			 | (OP==`LDA_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDA_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`LDA_aby & T==`Tfour & phi1)
			 | (OP==`LDY_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDY_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`LDY_abx & T==`Tfour & phi1)
			 | (OP==`LDA_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDA_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`LDA_abx & T==`Tfour & phi1)
			 | (OP==`LDX_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDX_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`LDX_aby & T==`Tfour & phi1)
			 | (OP==`CMP_izx & T==`Tzero & phi1)
			 | (OP==`CMP_izx & T==`Tthree & phi1)
			 | (OP==`CMP_izx & T==`Tfour & phi1)
			 | (OP==`CMP_izx & T==`Tfive & phi1)
			 | (OP==`CPY_zp & T==`Tzero & phi1)
			 | (OP==`CMP_zp & T==`Tzero & phi1)
			 | (OP==`DEC_zp & T==`Tzero & phi1)
			 | (OP==`DEC_zp & T==`Tthree & phi1)
			 | (OP==`DEC_zp & T==`Tfour & phi1)
			 | (OP==`CPY_abs & T==`Tzero & phi1)
			 | (OP==`CMP_abs & T==`Tzero & phi1)
			 | (OP==`DEC_abs & T==`Tzero & phi1)
			 | (OP==`DEC_abs & T==`Tfour & phi1)
			 | (OP==`DEC_abs & T==`Tfive & phi1)
			 | (OP==`CMP_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`CMP_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`CMP_izy & T==`Tthree & phi1)
			 | (OP==`CMP_izy & T==`Tfour & phi1)
			 | (OP==`CMP_izy & T==`Tfive & phi1)
			 | (OP==`CMP_zpx & T==`Tzero & phi1)
			 | (OP==`CMP_zpx & T==`Tthree & phi1)
			 | (OP==`DEC_zpx & T==`Tzero & phi1)
			 | (OP==`DEC_zpx & T==`Tthree & phi1)
			 | (OP==`DEC_zpx & T==`Tfour & phi1)
			 | (OP==`DEC_zpx & T==`Tfive & phi1)
			 | (OP==`CMP_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`CMP_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`CMP_aby & T==`Tfour & phi1)
			 | (OP==`CMP_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`CMP_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`CMP_abx & T==`Tfour & phi1)
			 | (OP==`DEC_abx & T==`Tzero & phi1)
			 | (OP==`DEC_abx & T==`Tfour & phi1)
			 | (OP==`DEC_abx & T==`Tfive & phi1)
			 | (OP==`DEC_abx & T==`Tsix & phi1)
			 | (OP==`SBC_izx & T==`Tzero & phi1)
			 | (OP==`SBC_izx & T==`Tthree & phi1)
			 | (OP==`SBC_izx & T==`Tfour & phi1)
			 | (OP==`SBC_izx & T==`Tfive & phi1)
			 | (OP==`CPX_zp & T==`Tzero & phi1)
			 | (OP==`SBC_zp & T==`Tzero & phi1)
			 | (OP==`INC_zp & T==`Tzero & phi1)
			 | (OP==`INC_zp & T==`Tthree & phi1)
			 | (OP==`INC_zp & T==`Tfour & phi1)
			 | (OP==`CPX_abs & T==`Tzero & phi1)
			 | (OP==`SBC_abs & T==`Tzero & phi1)
			 | (OP==`INC_abs & T==`Tzero & phi1)
			 | (OP==`INC_abs & T==`Tfour & phi1)
			 | (OP==`INC_abs & T==`Tfive & phi1)
			 | (OP==`SBC_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`SBC_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`SBC_izy & T==`Tthree & phi1)
			 | (OP==`SBC_izy & T==`Tfour & phi1)
			 | (OP==`SBC_izy & T==`Tfive & phi1)
			 | (OP==`SBC_zpx & T==`Tzero & phi1)
			 | (OP==`SBC_zpx & T==`Tthree & phi1)
			 | (OP==`INC_zpx & T==`Tzero & phi1)
			 | (OP==`INC_zpx & T==`Tthree & phi1)
			 | (OP==`INC_zpx & T==`Tfour & phi1)
			 | (OP==`INC_zpx & T==`Tfive & phi1)
			 | (OP==`SBC_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`SBC_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`SBC_aby & T==`Tfour & phi1)
			 | (OP==`SBC_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`SBC_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`SBC_abx & T==`Tfour & phi1)
			 | (OP==`INC_abx & T==`Tzero & phi1)
			 | (OP==`INC_abx & T==`Tfour & phi1)
			 | (OP==`INC_abx & T==`Tfive & phi1)
			 | (OP==`INC_abx & T==`Tsix & phi1)
			;

assign control[`ADL_PCL] = (OP==`BRK & T==`Tone & phi1)
			 | (OP==`BRK & T==`Ttwo & phi1)
			 | (OP==`ORA_izx & T==`Tone & phi1)
			 | (OP==`ORA_izx & T==`Ttwo & phi1)
			 | (OP==`ORA_zp & T==`Tone & phi1)
			 | (OP==`ORA_zp & T==`Ttwo & phi1)
			 | (OP==`ASL_zp & T==`Tone & phi1)
			 | (OP==`ASL_zp & T==`Ttwo & phi1)
			 | (OP==`PHP & T==`Tone & phi1)
			 | (OP==`PHP & T==`Ttwo & phi1)
			 | (OP==`ORA_imm & T==`Tone & phi1)
			 | (OP==`ORA_imm & T==`Ttwo & phi1)
			 | (OP==`ASL & T==`Tone & phi1)
			 | (OP==`ASL & T==`Ttwo & phi1)
			 | (OP==`ORA_abs & T==`Tone & phi1)
			 | (OP==`ORA_abs & T==`Ttwo & phi1)
			 | (OP==`ORA_abs & T==`Tthree & phi1)
			 | (OP==`ASL_abs & T==`Tone & phi1)
			 | (OP==`ASL_abs & T==`Ttwo & phi1)
			 | (OP==`ASL_abs & T==`Tthree & phi1)
			 | (OP==`BPL_rel & T==`Tzero & phi1)
			 | (OP==`BPL_rel & T==`Ttwo & phi1)
			 | (OP==`BPL_rel & T==`Tthree & phi1)
			 | (OP==`BPL_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BPL_rel & T==`T1BranchCross & phi1)
			 | (OP==`BPL_rel & T==`T1NoBranch & phi1)
			 | (OP==`ORA_izy & T==`Tone & phi1)
			 | (OP==`ORA_izy & T==`Ttwo & phi1)
			 | (OP==`ORA_zpx & T==`Tone & phi1)
			 | (OP==`ORA_zpx & T==`Ttwo & phi1)
			 | (OP==`ASL_zpx & T==`Tone & phi1)
			 | (OP==`ASL_zpx & T==`Ttwo & phi1)
			 | (OP==`CLC & T==`Tone & phi1)
			 | (OP==`CLC & T==`Ttwo & phi1)
			 | (OP==`ORA_aby & T==`Tone & phi1)
			 | (OP==`ORA_aby & T==`Ttwo & phi1)
			 | (OP==`ORA_aby & T==`Tthree & phi1)
			 | (OP==`ORA_abx & T==`Tone & phi1)
			 | (OP==`ORA_abx & T==`Ttwo & phi1)
			 | (OP==`ORA_abx & T==`Tthree & phi1)
			 | (OP==`ASL_abx & T==`Tone & phi1)
			 | (OP==`ASL_abx & T==`Ttwo & phi1)
			 | (OP==`ASL_abx & T==`Tthree & phi1)
			 | (OP==`JSR_abs & T==`Tzero & phi1)
			 | (OP==`JSR_abs & T==`Tone & phi1)
			 | (OP==`JSR_abs & T==`Ttwo & phi1)
			 | (OP==`AND_izx & T==`Tone & phi1)
			 | (OP==`AND_izx & T==`Ttwo & phi1)
			 | (OP==`BIT_zp & T==`Tone & phi1)
			 | (OP==`BIT_zp & T==`Ttwo & phi1)
			 | (OP==`AND_zp & T==`Tone & phi1)
			 | (OP==`AND_zp & T==`Ttwo & phi1)
			 | (OP==`ROL_zp & T==`Tone & phi1)
			 | (OP==`ROL_zp & T==`Ttwo & phi1)
			 | (OP==`PLP & T==`Tone & phi1)
			 | (OP==`PLP & T==`Ttwo & phi1)
			 | (OP==`AND_imm & T==`Tone & phi1)
			 | (OP==`AND_imm & T==`Ttwo & phi1)
			 | (OP==`ROL & T==`Tone & phi1)
			 | (OP==`ROL & T==`Ttwo & phi1)
			 | (OP==`BIT_abs & T==`Tone & phi1)
			 | (OP==`BIT_abs & T==`Ttwo & phi1)
			 | (OP==`BIT_abs & T==`Tthree & phi1)
			 | (OP==`AND_abs & T==`Tone & phi1)
			 | (OP==`AND_abs & T==`Ttwo & phi1)
			 | (OP==`AND_abs & T==`Tthree & phi1)
			 | (OP==`ROL_abs & T==`Tone & phi1)
			 | (OP==`ROL_abs & T==`Ttwo & phi1)
			 | (OP==`ROL_abs & T==`Tthree & phi1)
			 | (OP==`BMI_rel & T==`Tzero & phi1)
			 | (OP==`BMI_rel & T==`Ttwo & phi1)
			 | (OP==`BMI_rel & T==`Tthree & phi1)
			 | (OP==`BMI_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BMI_rel & T==`T1BranchCross & phi1)
			 | (OP==`BMI_rel & T==`T1NoBranch & phi1)
			 | (OP==`AND_izy & T==`Tone & phi1)
			 | (OP==`AND_izy & T==`Ttwo & phi1)
			 | (OP==`AND_zpx & T==`Tone & phi1)
			 | (OP==`AND_zpx & T==`Ttwo & phi1)
			 | (OP==`ROL_zpx & T==`Tone & phi1)
			 | (OP==`ROL_zpx & T==`Ttwo & phi1)
			 | (OP==`SEC & T==`Tone & phi1)
			 | (OP==`SEC & T==`Ttwo & phi1)
			 | (OP==`AND_aby & T==`Tone & phi1)
			 | (OP==`AND_aby & T==`Ttwo & phi1)
			 | (OP==`AND_aby & T==`Tthree & phi1)
			 | (OP==`AND_abx & T==`Tone & phi1)
			 | (OP==`AND_abx & T==`Ttwo & phi1)
			 | (OP==`AND_abx & T==`Tthree & phi1)
			 | (OP==`ROL_abx & T==`Tone & phi1)
			 | (OP==`ROL_abx & T==`Ttwo & phi1)
			 | (OP==`ROL_abx & T==`Tthree & phi1)
			 | (OP==`RTI & T==`Tone & phi1)
			 | (OP==`RTI & T==`Ttwo & phi1)
			 | (OP==`EOR_izx & T==`Tone & phi1)
			 | (OP==`EOR_izx & T==`Ttwo & phi1)
			 | (OP==`EOR_zp & T==`Tone & phi1)
			 | (OP==`EOR_zp & T==`Ttwo & phi1)
			 | (OP==`LSR_zp & T==`Tone & phi1)
			 | (OP==`LSR_zp & T==`Ttwo & phi1)
			 | (OP==`PHA & T==`Tone & phi1)
			 | (OP==`PHA & T==`Ttwo & phi1)
			 | (OP==`EOR_imm & T==`Tone & phi1)
			 | (OP==`EOR_imm & T==`Ttwo & phi1)
			 | (OP==`LSR & T==`Tone & phi1)
			 | (OP==`LSR & T==`Ttwo & phi1)
			 | (OP==`JMP_abs & T==`Tzero & phi1)
			 | (OP==`JMP_abs & T==`Tone & phi1)
			 | (OP==`JMP_abs & T==`Ttwo & phi1)
			 | (OP==`EOR_abs & T==`Tone & phi1)
			 | (OP==`EOR_abs & T==`Ttwo & phi1)
			 | (OP==`EOR_abs & T==`Tthree & phi1)
			 | (OP==`LSR_abs & T==`Tone & phi1)
			 | (OP==`LSR_abs & T==`Ttwo & phi1)
			 | (OP==`LSR_abs & T==`Tthree & phi1)
			 | (OP==`BVC_rel & T==`Tzero & phi1)
			 | (OP==`BVC_rel & T==`Ttwo & phi1)
			 | (OP==`BVC_rel & T==`Tthree & phi1)
			 | (OP==`BVC_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BVC_rel & T==`T1BranchCross & phi1)
			 | (OP==`BVC_rel & T==`T1NoBranch & phi1)
			 | (OP==`EOR_izy & T==`Tone & phi1)
			 | (OP==`EOR_izy & T==`Ttwo & phi1)
			 | (OP==`EOR_zpx & T==`Tone & phi1)
			 | (OP==`EOR_zpx & T==`Ttwo & phi1)
			 | (OP==`LSR_zpx & T==`Tone & phi1)
			 | (OP==`LSR_zpx & T==`Ttwo & phi1)
			 | (OP==`CLI & T==`Tone & phi1)
			 | (OP==`CLI & T==`Ttwo & phi1)
			 | (OP==`EOR_aby & T==`Tone & phi1)
			 | (OP==`EOR_aby & T==`Ttwo & phi1)
			 | (OP==`EOR_aby & T==`Tthree & phi1)
			 | (OP==`EOR_abx & T==`Tone & phi1)
			 | (OP==`EOR_abx & T==`Ttwo & phi1)
			 | (OP==`EOR_abx & T==`Tthree & phi1)
			 | (OP==`LSR_abx & T==`Tone & phi1)
			 | (OP==`LSR_abx & T==`Ttwo & phi1)
			 | (OP==`LSR_abx & T==`Tthree & phi1)
			 | (OP==`RTS & T==`Tzero & phi1)
			 | (OP==`RTS & T==`Tone & phi1)
			 | (OP==`RTS & T==`Ttwo & phi1)
			 | (OP==`ADC_izx & T==`Tone & phi1)
			 | (OP==`ADC_izx & T==`Ttwo & phi1)
			 | (OP==`ADC_zp & T==`Tone & phi1)
			 | (OP==`ADC_zp & T==`Ttwo & phi1)
			 | (OP==`ROR_zp & T==`Tone & phi1)
			 | (OP==`ROR_zp & T==`Ttwo & phi1)
			 | (OP==`PLA & T==`Tone & phi1)
			 | (OP==`PLA & T==`Ttwo & phi1)
			 | (OP==`ADC_imm & T==`Tone & phi1)
			 | (OP==`ADC_imm & T==`Ttwo & phi1)
			 | (OP==`ROR & T==`Tone & phi1)
			 | (OP==`ROR & T==`Ttwo & phi1)
			 | (OP==`JMP_zp & T==`Tone & phi1)
			 | (OP==`JMP_zp & T==`Ttwo & phi1)
			 | (OP==`JMP_zp & T==`Tthree & phi1)
			 | (OP==`ADC_abs & T==`Tone & phi1)
			 | (OP==`ADC_abs & T==`Ttwo & phi1)
			 | (OP==`ADC_abs & T==`Tthree & phi1)
			 | (OP==`ROR_abs & T==`Tone & phi1)
			 | (OP==`ROR_abs & T==`Ttwo & phi1)
			 | (OP==`ROR_abs & T==`Tthree & phi1)
			 | (OP==`BVS_rel & T==`Tzero & phi1)
			 | (OP==`BVS_rel & T==`Ttwo & phi1)
			 | (OP==`BVS_rel & T==`Tthree & phi1)
			 | (OP==`BVS_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BVS_rel & T==`T1BranchCross & phi1)
			 | (OP==`BVS_rel & T==`T1NoBranch & phi1)
			 | (OP==`ADC_izy & T==`Tone & phi1)
			 | (OP==`ADC_izy & T==`Ttwo & phi1)
			 | (OP==`ADC_zpx & T==`Tone & phi1)
			 | (OP==`ADC_zpx & T==`Ttwo & phi1)
			 | (OP==`ROR_zpx & T==`Tone & phi1)
			 | (OP==`ROR_zpx & T==`Ttwo & phi1)
			 | (OP==`SEI & T==`Tone & phi1)
			 | (OP==`SEI & T==`Ttwo & phi1)
			 | (OP==`ADC_aby & T==`Tone & phi1)
			 | (OP==`ADC_aby & T==`Ttwo & phi1)
			 | (OP==`ADC_aby & T==`Tthree & phi1)
			 | (OP==`ADC_abx & T==`Tone & phi1)
			 | (OP==`ADC_abx & T==`Ttwo & phi1)
			 | (OP==`ADC_abx & T==`Tthree & phi1)
			 | (OP==`ROR_abx & T==`Tone & phi1)
			 | (OP==`ROR_abx & T==`Ttwo & phi1)
			 | (OP==`ROR_abx & T==`Tthree & phi1)
			 | (OP==`STA_izx & T==`Tone & phi1)
			 | (OP==`STA_izx & T==`Ttwo & phi1)
			 | (OP==`STY_zp & T==`Tone & phi1)
			 | (OP==`STY_zp & T==`Ttwo & phi1)
			 | (OP==`STA_zp & T==`Tone & phi1)
			 | (OP==`STA_zp & T==`Ttwo & phi1)
			 | (OP==`STX_zp & T==`Tone & phi1)
			 | (OP==`STX_zp & T==`Ttwo & phi1)
			 | (OP==`DEY & T==`Tone & phi1)
			 | (OP==`DEY & T==`Ttwo & phi1)
			 | (OP==`TXA & T==`Tone & phi1)
			 | (OP==`TXA & T==`Ttwo & phi1)
			 | (OP==`STY_abs & T==`Tone & phi1)
			 | (OP==`STY_abs & T==`Ttwo & phi1)
			 | (OP==`STY_abs & T==`Tthree & phi1)
			 | (OP==`STA_abs & T==`Tone & phi1)
			 | (OP==`STA_abs & T==`Ttwo & phi1)
			 | (OP==`STA_abs & T==`Tthree & phi1)
			 | (OP==`STX_abs & T==`Tone & phi1)
			 | (OP==`STX_abs & T==`Ttwo & phi1)
			 | (OP==`STX_abs & T==`Tthree & phi1)
			 | (OP==`BCC_rel & T==`Tzero & phi1)
			 | (OP==`BCC_rel & T==`Ttwo & phi1)
			 | (OP==`BCC_rel & T==`Tthree & phi1)
			 | (OP==`BCC_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BCC_rel & T==`T1BranchCross & phi1)
			 | (OP==`BCC_rel & T==`T1NoBranch & phi1)
			 | (OP==`STA_izy & T==`Tone & phi1)
			 | (OP==`STA_izy & T==`Ttwo & phi1)
			 | (OP==`STY_zpx & T==`Tone & phi1)
			 | (OP==`STY_zpx & T==`Ttwo & phi1)
			 | (OP==`STA_zpx & T==`Tone & phi1)
			 | (OP==`STA_zpx & T==`Ttwo & phi1)
			 | (OP==`STX_zpy & T==`Tone & phi1)
			 | (OP==`STX_zpy & T==`Ttwo & phi1)
			 | (OP==`TYA & T==`Tone & phi1)
			 | (OP==`TYA & T==`Ttwo & phi1)
			 | (OP==`STA_aby & T==`Tone & phi1)
			 | (OP==`STA_aby & T==`Ttwo & phi1)
			 | (OP==`STA_aby & T==`Tthree & phi1)
			 | (OP==`TXS & T==`Tone & phi1)
			 | (OP==`TXS & T==`Ttwo & phi1)
			 | (OP==`STA_abx & T==`Tone & phi1)
			 | (OP==`STA_abx & T==`Ttwo & phi1)
			 | (OP==`STA_abx & T==`Tthree & phi1)
			 | (OP==`LDY_imm & T==`Tone & phi1)
			 | (OP==`LDY_imm & T==`Ttwo & phi1)
			 | (OP==`LDA_izx & T==`Tone & phi1)
			 | (OP==`LDA_izx & T==`Ttwo & phi1)
			 | (OP==`LDX_imm & T==`Tone & phi1)
			 | (OP==`LDX_imm & T==`Ttwo & phi1)
			 | (OP==`LDY_zp & T==`Tone & phi1)
			 | (OP==`LDY_zp & T==`Ttwo & phi1)
			 | (OP==`LDA_zp & T==`Tone & phi1)
			 | (OP==`LDA_zp & T==`Ttwo & phi1)
			 | (OP==`LDX_zp & T==`Tone & phi1)
			 | (OP==`LDX_zp & T==`Ttwo & phi1)
			 | (OP==`TAY & T==`Tone & phi1)
			 | (OP==`TAY & T==`Ttwo & phi1)
			 | (OP==`LDA_imm & T==`Tone & phi1)
			 | (OP==`LDA_imm & T==`Ttwo & phi1)
			 | (OP==`TAX & T==`Tone & phi1)
			 | (OP==`TAX & T==`Ttwo & phi1)
			 | (OP==`LDY_abs & T==`Tone & phi1)
			 | (OP==`LDY_abs & T==`Ttwo & phi1)
			 | (OP==`LDY_abs & T==`Tthree & phi1)
			 | (OP==`LDA_abs & T==`Tone & phi1)
			 | (OP==`LDA_abs & T==`Ttwo & phi1)
			 | (OP==`LDA_abs & T==`Tthree & phi1)
			 | (OP==`LDX_abs & T==`Tone & phi1)
			 | (OP==`LDX_abs & T==`Ttwo & phi1)
			 | (OP==`LDX_abs & T==`Tthree & phi1)
			 | (OP==`BCS_rel & T==`Tzero & phi1)
			 | (OP==`BCS_rel & T==`Ttwo & phi1)
			 | (OP==`BCS_rel & T==`Tthree & phi1)
			 | (OP==`BCS_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BCS_rel & T==`T1BranchCross & phi1)
			 | (OP==`BCS_rel & T==`T1NoBranch & phi1)
			 | (OP==`LDA_izy & T==`Tone & phi1)
			 | (OP==`LDA_izy & T==`Ttwo & phi1)
			 | (OP==`LDY_zpx & T==`Tone & phi1)
			 | (OP==`LDY_zpx & T==`Ttwo & phi1)
			 | (OP==`LDA_zpx & T==`Tone & phi1)
			 | (OP==`LDA_zpx & T==`Ttwo & phi1)
			 | (OP==`LDX_zpy & T==`Tone & phi1)
			 | (OP==`LDX_zpy & T==`Ttwo & phi1)
			 | (OP==`CLV & T==`Tone & phi1)
			 | (OP==`CLV & T==`Ttwo & phi1)
			 | (OP==`LDA_aby & T==`Tone & phi1)
			 | (OP==`LDA_aby & T==`Ttwo & phi1)
			 | (OP==`LDA_aby & T==`Tthree & phi1)
			 | (OP==`TSX & T==`Tone & phi1)
			 | (OP==`TSX & T==`Ttwo & phi1)
			 | (OP==`LDY_abx & T==`Tone & phi1)
			 | (OP==`LDY_abx & T==`Ttwo & phi1)
			 | (OP==`LDY_abx & T==`Tthree & phi1)
			 | (OP==`LDA_abx & T==`Tone & phi1)
			 | (OP==`LDA_abx & T==`Ttwo & phi1)
			 | (OP==`LDA_abx & T==`Tthree & phi1)
			 | (OP==`LDX_aby & T==`Tone & phi1)
			 | (OP==`LDX_aby & T==`Ttwo & phi1)
			 | (OP==`LDX_aby & T==`Tthree & phi1)
			 | (OP==`CPY_imm & T==`Tone & phi1)
			 | (OP==`CPY_imm & T==`Ttwo & phi1)
			 | (OP==`CMP_izx & T==`Tone & phi1)
			 | (OP==`CMP_izx & T==`Ttwo & phi1)
			 | (OP==`CPY_zp & T==`Tone & phi1)
			 | (OP==`CPY_zp & T==`Ttwo & phi1)
			 | (OP==`CMP_zp & T==`Tone & phi1)
			 | (OP==`CMP_zp & T==`Ttwo & phi1)
			 | (OP==`DEC_zp & T==`Tone & phi1)
			 | (OP==`DEC_zp & T==`Ttwo & phi1)
			 | (OP==`INY & T==`Tone & phi1)
			 | (OP==`INY & T==`Ttwo & phi1)
			 | (OP==`CMP_imm & T==`Tone & phi1)
			 | (OP==`CMP_imm & T==`Ttwo & phi1)
			 | (OP==`DEX & T==`Tone & phi1)
			 | (OP==`DEX & T==`Ttwo & phi1)
			 | (OP==`CPY_abs & T==`Tone & phi1)
			 | (OP==`CPY_abs & T==`Ttwo & phi1)
			 | (OP==`CPY_abs & T==`Tthree & phi1)
			 | (OP==`CMP_abs & T==`Tone & phi1)
			 | (OP==`CMP_abs & T==`Ttwo & phi1)
			 | (OP==`CMP_abs & T==`Tthree & phi1)
			 | (OP==`DEC_abs & T==`Tone & phi1)
			 | (OP==`DEC_abs & T==`Ttwo & phi1)
			 | (OP==`DEC_abs & T==`Tthree & phi1)
			 | (OP==`BNE_rel & T==`Tzero & phi1)
			 | (OP==`BNE_rel & T==`Ttwo & phi1)
			 | (OP==`BNE_rel & T==`Tthree & phi1)
			 | (OP==`BNE_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BNE_rel & T==`T1BranchCross & phi1)
			 | (OP==`BNE_rel & T==`T1NoBranch & phi1)
			 | (OP==`CMP_izy & T==`Tone & phi1)
			 | (OP==`CMP_izy & T==`Ttwo & phi1)
			 | (OP==`CMP_zpx & T==`Tone & phi1)
			 | (OP==`CMP_zpx & T==`Ttwo & phi1)
			 | (OP==`DEC_zpx & T==`Tone & phi1)
			 | (OP==`DEC_zpx & T==`Ttwo & phi1)
			 | (OP==`CLD & T==`Tone & phi1)
			 | (OP==`CLD & T==`Ttwo & phi1)
			 | (OP==`CMP_aby & T==`Tone & phi1)
			 | (OP==`CMP_aby & T==`Ttwo & phi1)
			 | (OP==`CMP_aby & T==`Tthree & phi1)
			 | (OP==`CMP_abx & T==`Tone & phi1)
			 | (OP==`CMP_abx & T==`Ttwo & phi1)
			 | (OP==`CMP_abx & T==`Tthree & phi1)
			 | (OP==`DEC_abx & T==`Tone & phi1)
			 | (OP==`DEC_abx & T==`Ttwo & phi1)
			 | (OP==`DEC_abx & T==`Tthree & phi1)
			 | (OP==`CPX_imm & T==`Tone & phi1)
			 | (OP==`CPX_imm & T==`Ttwo & phi1)
			 | (OP==`SBC_izx & T==`Tone & phi1)
			 | (OP==`SBC_izx & T==`Ttwo & phi1)
			 | (OP==`CPX_zp & T==`Tone & phi1)
			 | (OP==`CPX_zp & T==`Ttwo & phi1)
			 | (OP==`SBC_zp & T==`Tone & phi1)
			 | (OP==`SBC_zp & T==`Ttwo & phi1)
			 | (OP==`INC_zp & T==`Tone & phi1)
			 | (OP==`INC_zp & T==`Ttwo & phi1)
			 | (OP==`INX & T==`Tone & phi1)
			 | (OP==`INX & T==`Ttwo & phi1)
			 | (OP==`SBC_imm & T==`Tone & phi1)
			 | (OP==`SBC_imm & T==`Ttwo & phi1)
			 | (OP==`NOP & T==`Tone & phi1)
			 | (OP==`NOP & T==`Ttwo & phi1)
			 | (OP==`CPX_abs & T==`Tone & phi1)
			 | (OP==`CPX_abs & T==`Ttwo & phi1)
			 | (OP==`CPX_abs & T==`Tthree & phi1)
			 | (OP==`SBC_abs & T==`Tone & phi1)
			 | (OP==`SBC_abs & T==`Ttwo & phi1)
			 | (OP==`SBC_abs & T==`Tthree & phi1)
			 | (OP==`INC_abs & T==`Tone & phi1)
			 | (OP==`INC_abs & T==`Ttwo & phi1)
			 | (OP==`INC_abs & T==`Tthree & phi1)
			 | (OP==`BEQ_rel & T==`Tzero & phi1)
			 | (OP==`BEQ_rel & T==`Ttwo & phi1)
			 | (OP==`BEQ_rel & T==`Tthree & phi1)
			 | (OP==`BEQ_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BEQ_rel & T==`T1BranchCross & phi1)
			 | (OP==`BEQ_rel & T==`T1NoBranch & phi1)
			 | (OP==`SBC_izy & T==`Tone & phi1)
			 | (OP==`SBC_izy & T==`Ttwo & phi1)
			 | (OP==`SBC_zpx & T==`Tone & phi1)
			 | (OP==`SBC_zpx & T==`Ttwo & phi1)
			 | (OP==`INC_zpx & T==`Tone & phi1)
			 | (OP==`INC_zpx & T==`Ttwo & phi1)
			 | (OP==`SED & T==`Tone & phi1)
			 | (OP==`SED & T==`Ttwo & phi1)
			 | (OP==`SBC_aby & T==`Tone & phi1)
			 | (OP==`SBC_aby & T==`Ttwo & phi1)
			 | (OP==`SBC_aby & T==`Tthree & phi1)
			 | (OP==`SBC_abx & T==`Tone & phi1)
			 | (OP==`SBC_abx & T==`Ttwo & phi1)
			 | (OP==`SBC_abx & T==`Tthree & phi1)
			 | (OP==`INC_abx & T==`Tone & phi1)
			 | (OP==`INC_abx & T==`Ttwo & phi1)
			 | (OP==`INC_abx & T==`Tthree & phi1)
			;

assign control[`nI_PC] = (OP==`BRK & T==`Tzero & phi1)
			 | (OP==`BRK & T==`Tzero & phi2)
			 | (OP==`BRK & T==`Tthree & phi1)
			 | (OP==`BRK & T==`Tthree & phi2)
			 | (OP==`BRK & T==`Tfour & phi1)
			 | (OP==`BRK & T==`Tfour & phi2)
			 | (OP==`BRK & T==`Tfive & phi1)
			 | (OP==`BRK & T==`Tfive & phi2)
			 | (OP==`BRK & T==`Tsix & phi1)
			 | (OP==`BRK & T==`Tsix & phi2)
			 | (OP==`ORA_izx & T==`Tzero & phi1)
			 | (OP==`ORA_izx & T==`Tzero & phi2)
			 | (OP==`ORA_izx & T==`Tthree & phi1)
			 | (OP==`ORA_izx & T==`Tthree & phi2)
			 | (OP==`ORA_izx & T==`Tfour & phi1)
			 | (OP==`ORA_izx & T==`Tfour & phi2)
			 | (OP==`ORA_izx & T==`Tfive & phi1)
			 | (OP==`ORA_izx & T==`Tfive & phi2)
			 | (OP==`ORA_zp & T==`Tzero & phi1)
			 | (OP==`ORA_zp & T==`Tzero & phi2)
			 | (OP==`ASL_zp & T==`Tzero & phi1)
			 | (OP==`ASL_zp & T==`Tzero & phi2)
			 | (OP==`ASL_zp & T==`Tthree & phi1)
			 | (OP==`ASL_zp & T==`Tthree & phi2)
			 | (OP==`ASL_zp & T==`Tfour & phi1)
			 | (OP==`ASL_zp & T==`Tfour & phi2)
			 | (OP==`PHP & T==`Tzero & phi1)
			 | (OP==`PHP & T==`Tzero & phi2)
			 | (OP==`PHP & T==`Ttwo & phi1)
			 | (OP==`PHP & T==`Ttwo & phi2)
			 | (OP==`ASL & T==`Ttwo & phi1)
			 | (OP==`ASL & T==`Ttwo & phi2)
			 | (OP==`ORA_abs & T==`Tzero & phi1)
			 | (OP==`ORA_abs & T==`Tzero & phi2)
			 | (OP==`ASL_abs & T==`Tzero & phi1)
			 | (OP==`ASL_abs & T==`Tzero & phi2)
			 | (OP==`ASL_abs & T==`Tfour & phi1)
			 | (OP==`ASL_abs & T==`Tfour & phi2)
			 | (OP==`ASL_abs & T==`Tfive & phi1)
			 | (OP==`ASL_abs & T==`Tfive & phi2)
			 | (OP==`BPL_rel & T==`Tzero & phi1)
			 | (OP==`BPL_rel & T==`Tzero & phi2)
			 | (OP==`BPL_rel & T==`Tthree & phi1)
			 | (OP==`BPL_rel & T==`Tthree & phi2)
			 | (OP==`ORA_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`ORA_izy & T==`TzeroCrossPg & phi2)
			 | (OP==`ORA_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ORA_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`ORA_izy & T==`Tthree & phi1)
			 | (OP==`ORA_izy & T==`Tthree & phi2)
			 | (OP==`ORA_izy & T==`Tfour & phi1)
			 | (OP==`ORA_izy & T==`Tfour & phi2)
			 | (OP==`ORA_izy & T==`Tfive & phi1)
			 | (OP==`ORA_izy & T==`Tfive & phi2)
			 | (OP==`ORA_zpx & T==`Tzero & phi1)
			 | (OP==`ORA_zpx & T==`Tzero & phi2)
			 | (OP==`ORA_zpx & T==`Tthree & phi1)
			 | (OP==`ORA_zpx & T==`Tthree & phi2)
			 | (OP==`ASL_zpx & T==`Tzero & phi1)
			 | (OP==`ASL_zpx & T==`Tzero & phi2)
			 | (OP==`ASL_zpx & T==`Tthree & phi1)
			 | (OP==`ASL_zpx & T==`Tthree & phi2)
			 | (OP==`ASL_zpx & T==`Tfour & phi1)
			 | (OP==`ASL_zpx & T==`Tfour & phi2)
			 | (OP==`ASL_zpx & T==`Tfive & phi1)
			 | (OP==`ASL_zpx & T==`Tfive & phi2)
			 | (OP==`CLC & T==`Ttwo & phi1)
			 | (OP==`CLC & T==`Ttwo & phi2)
			 | (OP==`ORA_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ORA_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`ORA_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`ORA_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`ORA_aby & T==`Tfour & phi1)
			 | (OP==`ORA_aby & T==`Tfour & phi2)
			 | (OP==`ORA_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ORA_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`ORA_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`ORA_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`ORA_abx & T==`Tfour & phi1)
			 | (OP==`ORA_abx & T==`Tfour & phi2)
			 | (OP==`ASL_abx & T==`Tzero & phi1)
			 | (OP==`ASL_abx & T==`Tzero & phi2)
			 | (OP==`ASL_abx & T==`Tfour & phi1)
			 | (OP==`ASL_abx & T==`Tfour & phi2)
			 | (OP==`ASL_abx & T==`Tfive & phi1)
			 | (OP==`ASL_abx & T==`Tfive & phi2)
			 | (OP==`ASL_abx & T==`Tsix & phi1)
			 | (OP==`ASL_abx & T==`Tsix & phi2)
			 | (OP==`JSR_abs & T==`Tthree & phi1)
			 | (OP==`JSR_abs & T==`Tthree & phi2)
			 | (OP==`JSR_abs & T==`Tfour & phi1)
			 | (OP==`JSR_abs & T==`Tfour & phi2)
			 | (OP==`JSR_abs & T==`Tfive & phi1)
			 | (OP==`JSR_abs & T==`Tfive & phi2)
			 | (OP==`AND_izx & T==`Tzero & phi1)
			 | (OP==`AND_izx & T==`Tzero & phi2)
			 | (OP==`AND_izx & T==`Tthree & phi1)
			 | (OP==`AND_izx & T==`Tthree & phi2)
			 | (OP==`AND_izx & T==`Tfour & phi1)
			 | (OP==`AND_izx & T==`Tfour & phi2)
			 | (OP==`AND_izx & T==`Tfive & phi1)
			 | (OP==`AND_izx & T==`Tfive & phi2)
			 | (OP==`BIT_zp & T==`Tzero & phi1)
			 | (OP==`BIT_zp & T==`Tzero & phi2)
			 | (OP==`AND_zp & T==`Tzero & phi1)
			 | (OP==`AND_zp & T==`Tzero & phi2)
			 | (OP==`ROL_zp & T==`Tzero & phi1)
			 | (OP==`ROL_zp & T==`Tzero & phi2)
			 | (OP==`ROL_zp & T==`Tthree & phi1)
			 | (OP==`ROL_zp & T==`Tthree & phi2)
			 | (OP==`ROL_zp & T==`Tfour & phi1)
			 | (OP==`ROL_zp & T==`Tfour & phi2)
			 | (OP==`PLP & T==`Tzero & phi1)
			 | (OP==`PLP & T==`Tzero & phi2)
			 | (OP==`PLP & T==`Ttwo & phi1)
			 | (OP==`PLP & T==`Ttwo & phi2)
			 | (OP==`PLP & T==`Tthree & phi1)
			 | (OP==`PLP & T==`Tthree & phi2)
			 | (OP==`ROL & T==`Ttwo & phi1)
			 | (OP==`ROL & T==`Ttwo & phi2)
			 | (OP==`BIT_abs & T==`Tzero & phi1)
			 | (OP==`BIT_abs & T==`Tzero & phi2)
			 | (OP==`AND_abs & T==`Tzero & phi1)
			 | (OP==`AND_abs & T==`Tzero & phi2)
			 | (OP==`ROL_abs & T==`Tzero & phi1)
			 | (OP==`ROL_abs & T==`Tzero & phi2)
			 | (OP==`ROL_abs & T==`Tfour & phi1)
			 | (OP==`ROL_abs & T==`Tfour & phi2)
			 | (OP==`ROL_abs & T==`Tfive & phi1)
			 | (OP==`ROL_abs & T==`Tfive & phi2)
			 | (OP==`BMI_rel & T==`Tzero & phi1)
			 | (OP==`BMI_rel & T==`Tzero & phi2)
			 | (OP==`BMI_rel & T==`Tthree & phi1)
			 | (OP==`BMI_rel & T==`Tthree & phi2)
			 | (OP==`AND_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`AND_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`AND_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`AND_izy & T==`TzeroCrossPg & phi2)
			 | (OP==`AND_izy & T==`Tthree & phi1)
			 | (OP==`AND_izy & T==`Tthree & phi2)
			 | (OP==`AND_izy & T==`Tfour & phi1)
			 | (OP==`AND_izy & T==`Tfour & phi2)
			 | (OP==`AND_izy & T==`Tfive & phi1)
			 | (OP==`AND_izy & T==`Tfive & phi2)
			 | (OP==`AND_zpx & T==`Tzero & phi1)
			 | (OP==`AND_zpx & T==`Tzero & phi2)
			 | (OP==`AND_zpx & T==`Tthree & phi1)
			 | (OP==`AND_zpx & T==`Tthree & phi2)
			 | (OP==`ROL_zpx & T==`Tzero & phi1)
			 | (OP==`ROL_zpx & T==`Tzero & phi2)
			 | (OP==`ROL_zpx & T==`Tthree & phi1)
			 | (OP==`ROL_zpx & T==`Tthree & phi2)
			 | (OP==`ROL_zpx & T==`Tfour & phi1)
			 | (OP==`ROL_zpx & T==`Tfour & phi2)
			 | (OP==`ROL_zpx & T==`Tfive & phi1)
			 | (OP==`ROL_zpx & T==`Tfive & phi2)
			 | (OP==`SEC & T==`Ttwo & phi1)
			 | (OP==`SEC & T==`Ttwo & phi2)
			 | (OP==`AND_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`AND_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`AND_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`AND_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`AND_aby & T==`Tfour & phi1)
			 | (OP==`AND_aby & T==`Tfour & phi2)
			 | (OP==`AND_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`AND_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`AND_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`AND_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`AND_abx & T==`Tfour & phi1)
			 | (OP==`AND_abx & T==`Tfour & phi2)
			 | (OP==`ROL_abx & T==`Tzero & phi1)
			 | (OP==`ROL_abx & T==`Tzero & phi2)
			 | (OP==`ROL_abx & T==`Tfour & phi1)
			 | (OP==`ROL_abx & T==`Tfour & phi2)
			 | (OP==`ROL_abx & T==`Tfive & phi1)
			 | (OP==`ROL_abx & T==`Tfive & phi2)
			 | (OP==`ROL_abx & T==`Tsix & phi1)
			 | (OP==`ROL_abx & T==`Tsix & phi2)
			 | (OP==`RTI & T==`Tzero & phi1)
			 | (OP==`RTI & T==`Tzero & phi2)
			 | (OP==`RTI & T==`Tthree & phi1)
			 | (OP==`RTI & T==`Tthree & phi2)
			 | (OP==`RTI & T==`Tfour & phi1)
			 | (OP==`RTI & T==`Tfour & phi2)
			 | (OP==`RTI & T==`Tfive & phi1)
			 | (OP==`RTI & T==`Tfive & phi2)
			 | (OP==`EOR_izx & T==`Tzero & phi1)
			 | (OP==`EOR_izx & T==`Tzero & phi2)
			 | (OP==`EOR_izx & T==`Tthree & phi1)
			 | (OP==`EOR_izx & T==`Tthree & phi2)
			 | (OP==`EOR_izx & T==`Tfour & phi1)
			 | (OP==`EOR_izx & T==`Tfour & phi2)
			 | (OP==`EOR_izx & T==`Tfive & phi1)
			 | (OP==`EOR_izx & T==`Tfive & phi2)
			 | (OP==`EOR_zp & T==`Tzero & phi1)
			 | (OP==`EOR_zp & T==`Tzero & phi2)
			 | (OP==`LSR_zp & T==`Tzero & phi1)
			 | (OP==`LSR_zp & T==`Tzero & phi2)
			 | (OP==`LSR_zp & T==`Tthree & phi1)
			 | (OP==`LSR_zp & T==`Tthree & phi2)
			 | (OP==`LSR_zp & T==`Tfour & phi1)
			 | (OP==`LSR_zp & T==`Tfour & phi2)
			 | (OP==`PHA & T==`Tzero & phi1)
			 | (OP==`PHA & T==`Tzero & phi2)
			 | (OP==`PHA & T==`Ttwo & phi1)
			 | (OP==`PHA & T==`Ttwo & phi2)
			 | (OP==`LSR & T==`Ttwo & phi1)
			 | (OP==`LSR & T==`Ttwo & phi2)
			 | (OP==`EOR_abs & T==`Tzero & phi1)
			 | (OP==`EOR_abs & T==`Tzero & phi2)
			 | (OP==`LSR_abs & T==`Tzero & phi1)
			 | (OP==`LSR_abs & T==`Tzero & phi2)
			 | (OP==`LSR_abs & T==`Tfour & phi1)
			 | (OP==`LSR_abs & T==`Tfour & phi2)
			 | (OP==`LSR_abs & T==`Tfive & phi1)
			 | (OP==`LSR_abs & T==`Tfive & phi2)
			 | (OP==`BVC_rel & T==`Tzero & phi1)
			 | (OP==`BVC_rel & T==`Tzero & phi2)
			 | (OP==`BVC_rel & T==`Tthree & phi1)
			 | (OP==`BVC_rel & T==`Tthree & phi2)
			 | (OP==`EOR_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`EOR_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`EOR_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`EOR_izy & T==`TzeroCrossPg & phi2)
			 | (OP==`EOR_izy & T==`Tthree & phi1)
			 | (OP==`EOR_izy & T==`Tthree & phi2)
			 | (OP==`EOR_izy & T==`Tfour & phi1)
			 | (OP==`EOR_izy & T==`Tfour & phi2)
			 | (OP==`EOR_izy & T==`Tfive & phi1)
			 | (OP==`EOR_izy & T==`Tfive & phi2)
			 | (OP==`EOR_zpx & T==`Tzero & phi1)
			 | (OP==`EOR_zpx & T==`Tzero & phi2)
			 | (OP==`EOR_zpx & T==`Tthree & phi1)
			 | (OP==`EOR_zpx & T==`Tthree & phi2)
			 | (OP==`LSR_zpx & T==`Tzero & phi1)
			 | (OP==`LSR_zpx & T==`Tzero & phi2)
			 | (OP==`LSR_zpx & T==`Tthree & phi1)
			 | (OP==`LSR_zpx & T==`Tthree & phi2)
			 | (OP==`LSR_zpx & T==`Tfour & phi1)
			 | (OP==`LSR_zpx & T==`Tfour & phi2)
			 | (OP==`LSR_zpx & T==`Tfive & phi1)
			 | (OP==`LSR_zpx & T==`Tfive & phi2)
			 | (OP==`CLI & T==`Ttwo & phi1)
			 | (OP==`CLI & T==`Ttwo & phi2)
			 | (OP==`EOR_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`EOR_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`EOR_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`EOR_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`EOR_aby & T==`Tfour & phi1)
			 | (OP==`EOR_aby & T==`Tfour & phi2)
			 | (OP==`EOR_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`EOR_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`EOR_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`EOR_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`EOR_abx & T==`Tfour & phi1)
			 | (OP==`EOR_abx & T==`Tfour & phi2)
			 | (OP==`LSR_abx & T==`Tzero & phi1)
			 | (OP==`LSR_abx & T==`Tzero & phi2)
			 | (OP==`LSR_abx & T==`Tfour & phi1)
			 | (OP==`LSR_abx & T==`Tfour & phi2)
			 | (OP==`LSR_abx & T==`Tfive & phi1)
			 | (OP==`LSR_abx & T==`Tfive & phi2)
			 | (OP==`LSR_abx & T==`Tsix & phi1)
			 | (OP==`LSR_abx & T==`Tsix & phi2)
			 | (OP==`RTS & T==`Tthree & phi1)
			 | (OP==`RTS & T==`Tthree & phi2)
			 | (OP==`RTS & T==`Tfour & phi1)
			 | (OP==`RTS & T==`Tfour & phi2)
			 | (OP==`RTS & T==`Tfive & phi1)
			 | (OP==`RTS & T==`Tfive & phi2)
			 | (OP==`ADC_izx & T==`Tzero & phi1)
			 | (OP==`ADC_izx & T==`Tzero & phi2)
			 | (OP==`ADC_izx & T==`Tthree & phi1)
			 | (OP==`ADC_izx & T==`Tthree & phi2)
			 | (OP==`ADC_izx & T==`Tfour & phi1)
			 | (OP==`ADC_izx & T==`Tfour & phi2)
			 | (OP==`ADC_izx & T==`Tfive & phi1)
			 | (OP==`ADC_izx & T==`Tfive & phi2)
			 | (OP==`ADC_zp & T==`Tzero & phi1)
			 | (OP==`ADC_zp & T==`Tzero & phi2)
			 | (OP==`ROR_zp & T==`Tzero & phi1)
			 | (OP==`ROR_zp & T==`Tzero & phi2)
			 | (OP==`ROR_zp & T==`Tthree & phi1)
			 | (OP==`ROR_zp & T==`Tthree & phi2)
			 | (OP==`ROR_zp & T==`Tfour & phi1)
			 | (OP==`ROR_zp & T==`Tfour & phi2)
			 | (OP==`PLA & T==`Tzero & phi1)
			 | (OP==`PLA & T==`Tzero & phi2)
			 | (OP==`PLA & T==`Ttwo & phi1)
			 | (OP==`PLA & T==`Ttwo & phi2)
			 | (OP==`PLA & T==`Tthree & phi1)
			 | (OP==`PLA & T==`Tthree & phi2)
			 | (OP==`ROR & T==`Ttwo & phi1)
			 | (OP==`ROR & T==`Ttwo & phi2)
			 | (OP==`JMP_zp & T==`Tzero & phi1)
			 | (OP==`JMP_zp & T==`Tzero & phi2)
			 | (OP==`JMP_zp & T==`Tfour & phi1)
			 | (OP==`JMP_zp & T==`Tfour & phi2)
			 | (OP==`ADC_abs & T==`Tzero & phi1)
			 | (OP==`ADC_abs & T==`Tzero & phi2)
			 | (OP==`ROR_abs & T==`Tzero & phi1)
			 | (OP==`ROR_abs & T==`Tzero & phi2)
			 | (OP==`ROR_abs & T==`Tfour & phi1)
			 | (OP==`ROR_abs & T==`Tfour & phi2)
			 | (OP==`ROR_abs & T==`Tfive & phi1)
			 | (OP==`ROR_abs & T==`Tfive & phi2)
			 | (OP==`BVS_rel & T==`Tzero & phi1)
			 | (OP==`BVS_rel & T==`Tzero & phi2)
			 | (OP==`BVS_rel & T==`Tthree & phi1)
			 | (OP==`BVS_rel & T==`Tthree & phi2)
			 | (OP==`ADC_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ADC_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`ADC_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`ADC_izy & T==`TzeroCrossPg & phi2)
			 | (OP==`ADC_izy & T==`Tthree & phi1)
			 | (OP==`ADC_izy & T==`Tthree & phi2)
			 | (OP==`ADC_izy & T==`Tfour & phi1)
			 | (OP==`ADC_izy & T==`Tfour & phi2)
			 | (OP==`ADC_izy & T==`Tfive & phi1)
			 | (OP==`ADC_izy & T==`Tfive & phi2)
			 | (OP==`ADC_zpx & T==`Tzero & phi1)
			 | (OP==`ADC_zpx & T==`Tzero & phi2)
			 | (OP==`ADC_zpx & T==`Tthree & phi1)
			 | (OP==`ADC_zpx & T==`Tthree & phi2)
			 | (OP==`ROR_zpx & T==`Tzero & phi1)
			 | (OP==`ROR_zpx & T==`Tzero & phi2)
			 | (OP==`ROR_zpx & T==`Tthree & phi1)
			 | (OP==`ROR_zpx & T==`Tthree & phi2)
			 | (OP==`ROR_zpx & T==`Tfour & phi1)
			 | (OP==`ROR_zpx & T==`Tfour & phi2)
			 | (OP==`ROR_zpx & T==`Tfive & phi1)
			 | (OP==`ROR_zpx & T==`Tfive & phi2)
			 | (OP==`SEI & T==`Ttwo & phi1)
			 | (OP==`SEI & T==`Ttwo & phi2)
			 | (OP==`ADC_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ADC_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`ADC_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`ADC_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`ADC_aby & T==`Tfour & phi1)
			 | (OP==`ADC_aby & T==`Tfour & phi2)
			 | (OP==`ADC_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ADC_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`ADC_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`ADC_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`ADC_abx & T==`Tfour & phi1)
			 | (OP==`ADC_abx & T==`Tfour & phi2)
			 | (OP==`ROR_abx & T==`Tzero & phi1)
			 | (OP==`ROR_abx & T==`Tzero & phi2)
			 | (OP==`ROR_abx & T==`Tfour & phi1)
			 | (OP==`ROR_abx & T==`Tfour & phi2)
			 | (OP==`ROR_abx & T==`Tfive & phi1)
			 | (OP==`ROR_abx & T==`Tfive & phi2)
			 | (OP==`ROR_abx & T==`Tsix & phi1)
			 | (OP==`ROR_abx & T==`Tsix & phi2)
			 | (OP==`STA_izx & T==`Tzero & phi1)
			 | (OP==`STA_izx & T==`Tzero & phi2)
			 | (OP==`STA_izx & T==`Tthree & phi1)
			 | (OP==`STA_izx & T==`Tthree & phi2)
			 | (OP==`STA_izx & T==`Tfour & phi1)
			 | (OP==`STA_izx & T==`Tfour & phi2)
			 | (OP==`STA_izx & T==`Tfive & phi1)
			 | (OP==`STA_izx & T==`Tfive & phi2)
			 | (OP==`STY_zp & T==`Tzero & phi1)
			 | (OP==`STY_zp & T==`Tzero & phi2)
			 | (OP==`STA_zp & T==`Tzero & phi1)
			 | (OP==`STA_zp & T==`Tzero & phi2)
			 | (OP==`STX_zp & T==`Tzero & phi1)
			 | (OP==`STX_zp & T==`Tzero & phi2)
			 | (OP==`DEY & T==`Ttwo & phi1)
			 | (OP==`DEY & T==`Ttwo & phi2)
			 | (OP==`TXA & T==`Ttwo & phi1)
			 | (OP==`TXA & T==`Ttwo & phi2)
			 | (OP==`STY_abs & T==`Tzero & phi1)
			 | (OP==`STY_abs & T==`Tzero & phi2)
			 | (OP==`STA_abs & T==`Tzero & phi1)
			 | (OP==`STA_abs & T==`Tzero & phi2)
			 | (OP==`STX_abs & T==`Tzero & phi1)
			 | (OP==`STX_abs & T==`Tzero & phi2)
			 | (OP==`BCC_rel & T==`Tzero & phi1)
			 | (OP==`BCC_rel & T==`Tzero & phi2)
			 | (OP==`BCC_rel & T==`Tthree & phi1)
			 | (OP==`BCC_rel & T==`Tthree & phi2)
			 | (OP==`STA_izy & T==`Tzero & phi1)
			 | (OP==`STA_izy & T==`Tzero & phi2)
			 | (OP==`STA_izy & T==`Tthree & phi1)
			 | (OP==`STA_izy & T==`Tthree & phi2)
			 | (OP==`STA_izy & T==`Tfour & phi1)
			 | (OP==`STA_izy & T==`Tfour & phi2)
			 | (OP==`STA_izy & T==`Tfive & phi1)
			 | (OP==`STA_izy & T==`Tfive & phi2)
			 | (OP==`STY_zpx & T==`Tzero & phi1)
			 | (OP==`STY_zpx & T==`Tzero & phi2)
			 | (OP==`STY_zpx & T==`Tthree & phi1)
			 | (OP==`STY_zpx & T==`Tthree & phi2)
			 | (OP==`STA_zpx & T==`Tzero & phi1)
			 | (OP==`STA_zpx & T==`Tzero & phi2)
			 | (OP==`STA_zpx & T==`Tthree & phi1)
			 | (OP==`STA_zpx & T==`Tthree & phi2)
			 | (OP==`STX_zpy & T==`Tzero & phi1)
			 | (OP==`STX_zpy & T==`Tzero & phi2)
			 | (OP==`STX_zpy & T==`Tthree & phi1)
			 | (OP==`STX_zpy & T==`Tthree & phi2)
			 | (OP==`TYA & T==`Ttwo & phi1)
			 | (OP==`TYA & T==`Ttwo & phi2)
			 | (OP==`STA_aby & T==`Tzero & phi1)
			 | (OP==`STA_aby & T==`Tzero & phi2)
			 | (OP==`STA_aby & T==`Tfour & phi1)
			 | (OP==`STA_aby & T==`Tfour & phi2)
			 | (OP==`TXS & T==`Ttwo & phi1)
			 | (OP==`TXS & T==`Ttwo & phi2)
			 | (OP==`STA_abx & T==`Tzero & phi1)
			 | (OP==`STA_abx & T==`Tzero & phi2)
			 | (OP==`STA_abx & T==`Tfour & phi1)
			 | (OP==`STA_abx & T==`Tfour & phi2)
			 | (OP==`LDA_izx & T==`Tzero & phi1)
			 | (OP==`LDA_izx & T==`Tzero & phi2)
			 | (OP==`LDA_izx & T==`Tthree & phi1)
			 | (OP==`LDA_izx & T==`Tthree & phi2)
			 | (OP==`LDA_izx & T==`Tfour & phi1)
			 | (OP==`LDA_izx & T==`Tfour & phi2)
			 | (OP==`LDA_izx & T==`Tfive & phi1)
			 | (OP==`LDA_izx & T==`Tfive & phi2)
			 | (OP==`LDY_zp & T==`Tzero & phi1)
			 | (OP==`LDY_zp & T==`Tzero & phi2)
			 | (OP==`LDA_zp & T==`Tzero & phi1)
			 | (OP==`LDA_zp & T==`Tzero & phi2)
			 | (OP==`LDX_zp & T==`Tzero & phi1)
			 | (OP==`LDX_zp & T==`Tzero & phi2)
			 | (OP==`TAY & T==`Ttwo & phi1)
			 | (OP==`TAY & T==`Ttwo & phi2)
			 | (OP==`TAX & T==`Ttwo & phi1)
			 | (OP==`TAX & T==`Ttwo & phi2)
			 | (OP==`LDY_abs & T==`Tzero & phi1)
			 | (OP==`LDY_abs & T==`Tzero & phi2)
			 | (OP==`LDA_abs & T==`Tzero & phi1)
			 | (OP==`LDA_abs & T==`Tzero & phi2)
			 | (OP==`LDX_abs & T==`Tzero & phi1)
			 | (OP==`LDX_abs & T==`Tzero & phi2)
			 | (OP==`BCS_rel & T==`Tzero & phi1)
			 | (OP==`BCS_rel & T==`Tzero & phi2)
			 | (OP==`BCS_rel & T==`Tthree & phi1)
			 | (OP==`BCS_rel & T==`Tthree & phi2)
			 | (OP==`LDA_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDA_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`LDA_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`LDA_izy & T==`TzeroCrossPg & phi2)
			 | (OP==`LDA_izy & T==`Tthree & phi1)
			 | (OP==`LDA_izy & T==`Tthree & phi2)
			 | (OP==`LDA_izy & T==`Tfour & phi1)
			 | (OP==`LDA_izy & T==`Tfour & phi2)
			 | (OP==`LDA_izy & T==`Tfive & phi1)
			 | (OP==`LDA_izy & T==`Tfive & phi2)
			 | (OP==`LDY_zpx & T==`Tzero & phi1)
			 | (OP==`LDY_zpx & T==`Tzero & phi2)
			 | (OP==`LDY_zpx & T==`Tthree & phi1)
			 | (OP==`LDY_zpx & T==`Tthree & phi2)
			 | (OP==`LDA_zpx & T==`Tzero & phi1)
			 | (OP==`LDA_zpx & T==`Tzero & phi2)
			 | (OP==`LDA_zpx & T==`Tthree & phi1)
			 | (OP==`LDA_zpx & T==`Tthree & phi2)
			 | (OP==`LDX_zpy & T==`Tzero & phi1)
			 | (OP==`LDX_zpy & T==`Tzero & phi2)
			 | (OP==`LDX_zpy & T==`Tthree & phi1)
			 | (OP==`LDX_zpy & T==`Tthree & phi2)
			 | (OP==`CLV & T==`Ttwo & phi1)
			 | (OP==`CLV & T==`Ttwo & phi2)
			 | (OP==`LDA_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDA_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`LDA_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`LDA_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`LDA_aby & T==`Tfour & phi1)
			 | (OP==`LDA_aby & T==`Tfour & phi2)
			 | (OP==`TSX & T==`Ttwo & phi1)
			 | (OP==`TSX & T==`Ttwo & phi2)
			 | (OP==`LDY_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDY_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`LDY_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`LDY_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`LDY_abx & T==`Tfour & phi1)
			 | (OP==`LDY_abx & T==`Tfour & phi2)
			 | (OP==`LDA_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDA_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`LDA_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`LDA_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`LDA_abx & T==`Tfour & phi1)
			 | (OP==`LDA_abx & T==`Tfour & phi2)
			 | (OP==`LDX_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDX_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`LDX_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`LDX_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`LDX_aby & T==`Tfour & phi1)
			 | (OP==`LDX_aby & T==`Tfour & phi2)
			 | (OP==`CMP_izx & T==`Tzero & phi1)
			 | (OP==`CMP_izx & T==`Tzero & phi2)
			 | (OP==`CMP_izx & T==`Tthree & phi1)
			 | (OP==`CMP_izx & T==`Tthree & phi2)
			 | (OP==`CMP_izx & T==`Tfour & phi1)
			 | (OP==`CMP_izx & T==`Tfour & phi2)
			 | (OP==`CMP_izx & T==`Tfive & phi1)
			 | (OP==`CMP_izx & T==`Tfive & phi2)
			 | (OP==`CPY_zp & T==`Tzero & phi1)
			 | (OP==`CPY_zp & T==`Tzero & phi2)
			 | (OP==`CMP_zp & T==`Tzero & phi1)
			 | (OP==`CMP_zp & T==`Tzero & phi2)
			 | (OP==`DEC_zp & T==`Tzero & phi1)
			 | (OP==`DEC_zp & T==`Tzero & phi2)
			 | (OP==`DEC_zp & T==`Tthree & phi1)
			 | (OP==`DEC_zp & T==`Tthree & phi2)
			 | (OP==`DEC_zp & T==`Tfour & phi1)
			 | (OP==`DEC_zp & T==`Tfour & phi2)
			 | (OP==`INY & T==`Ttwo & phi1)
			 | (OP==`INY & T==`Ttwo & phi2)
			 | (OP==`DEX & T==`Ttwo & phi1)
			 | (OP==`DEX & T==`Ttwo & phi2)
			 | (OP==`CPY_abs & T==`Tzero & phi1)
			 | (OP==`CPY_abs & T==`Tzero & phi2)
			 | (OP==`CMP_abs & T==`Tzero & phi1)
			 | (OP==`CMP_abs & T==`Tzero & phi2)
			 | (OP==`DEC_abs & T==`Tzero & phi1)
			 | (OP==`DEC_abs & T==`Tzero & phi2)
			 | (OP==`DEC_abs & T==`Tfour & phi1)
			 | (OP==`DEC_abs & T==`Tfour & phi2)
			 | (OP==`DEC_abs & T==`Tfive & phi1)
			 | (OP==`DEC_abs & T==`Tfive & phi2)
			 | (OP==`BNE_rel & T==`Tzero & phi1)
			 | (OP==`BNE_rel & T==`Tzero & phi2)
			 | (OP==`BNE_rel & T==`Tthree & phi1)
			 | (OP==`BNE_rel & T==`Tthree & phi2)
			 | (OP==`CMP_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`CMP_izy & T==`TzeroCrossPg & phi2)
			 | (OP==`CMP_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`CMP_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`CMP_izy & T==`Tthree & phi1)
			 | (OP==`CMP_izy & T==`Tthree & phi2)
			 | (OP==`CMP_izy & T==`Tfour & phi1)
			 | (OP==`CMP_izy & T==`Tfour & phi2)
			 | (OP==`CMP_izy & T==`Tfive & phi1)
			 | (OP==`CMP_izy & T==`Tfive & phi2)
			 | (OP==`CMP_zpx & T==`Tzero & phi1)
			 | (OP==`CMP_zpx & T==`Tzero & phi2)
			 | (OP==`CMP_zpx & T==`Tthree & phi1)
			 | (OP==`CMP_zpx & T==`Tthree & phi2)
			 | (OP==`DEC_zpx & T==`Tzero & phi1)
			 | (OP==`DEC_zpx & T==`Tzero & phi2)
			 | (OP==`DEC_zpx & T==`Tthree & phi1)
			 | (OP==`DEC_zpx & T==`Tthree & phi2)
			 | (OP==`DEC_zpx & T==`Tfour & phi1)
			 | (OP==`DEC_zpx & T==`Tfour & phi2)
			 | (OP==`DEC_zpx & T==`Tfive & phi1)
			 | (OP==`DEC_zpx & T==`Tfive & phi2)
			 | (OP==`CLD & T==`Ttwo & phi1)
			 | (OP==`CLD & T==`Ttwo & phi2)
			 | (OP==`CMP_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`CMP_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`CMP_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`CMP_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`CMP_aby & T==`Tfour & phi1)
			 | (OP==`CMP_aby & T==`Tfour & phi2)
			 | (OP==`CMP_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`CMP_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`CMP_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`CMP_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`CMP_abx & T==`Tfour & phi1)
			 | (OP==`CMP_abx & T==`Tfour & phi2)
			 | (OP==`DEC_abx & T==`Tzero & phi1)
			 | (OP==`DEC_abx & T==`Tzero & phi2)
			 | (OP==`DEC_abx & T==`Tfour & phi1)
			 | (OP==`DEC_abx & T==`Tfour & phi2)
			 | (OP==`DEC_abx & T==`Tfive & phi1)
			 | (OP==`DEC_abx & T==`Tfive & phi2)
			 | (OP==`DEC_abx & T==`Tsix & phi1)
			 | (OP==`DEC_abx & T==`Tsix & phi2)
			 | (OP==`SBC_izx & T==`Tzero & phi1)
			 | (OP==`SBC_izx & T==`Tzero & phi2)
			 | (OP==`SBC_izx & T==`Tthree & phi1)
			 | (OP==`SBC_izx & T==`Tthree & phi2)
			 | (OP==`SBC_izx & T==`Tfour & phi1)
			 | (OP==`SBC_izx & T==`Tfour & phi2)
			 | (OP==`SBC_izx & T==`Tfive & phi1)
			 | (OP==`SBC_izx & T==`Tfive & phi2)
			 | (OP==`CPX_zp & T==`Tzero & phi1)
			 | (OP==`CPX_zp & T==`Tzero & phi2)
			 | (OP==`SBC_zp & T==`Tzero & phi1)
			 | (OP==`SBC_zp & T==`Tzero & phi2)
			 | (OP==`INC_zp & T==`Tzero & phi1)
			 | (OP==`INC_zp & T==`Tzero & phi2)
			 | (OP==`INC_zp & T==`Tthree & phi1)
			 | (OP==`INC_zp & T==`Tthree & phi2)
			 | (OP==`INC_zp & T==`Tfour & phi1)
			 | (OP==`INC_zp & T==`Tfour & phi2)
			 | (OP==`INX & T==`Ttwo & phi1)
			 | (OP==`INX & T==`Ttwo & phi2)
			 | (OP==`NOP & T==`Ttwo & phi1)
			 | (OP==`NOP & T==`Ttwo & phi2)
			 | (OP==`CPX_abs & T==`Tzero & phi1)
			 | (OP==`CPX_abs & T==`Tzero & phi2)
			 | (OP==`SBC_abs & T==`Tzero & phi1)
			 | (OP==`SBC_abs & T==`Tzero & phi2)
			 | (OP==`INC_abs & T==`Tzero & phi1)
			 | (OP==`INC_abs & T==`Tzero & phi2)
			 | (OP==`INC_abs & T==`Tfour & phi1)
			 | (OP==`INC_abs & T==`Tfour & phi2)
			 | (OP==`INC_abs & T==`Tfive & phi1)
			 | (OP==`INC_abs & T==`Tfive & phi2)
			 | (OP==`BEQ_rel & T==`Tzero & phi1)
			 | (OP==`BEQ_rel & T==`Tzero & phi2)
			 | (OP==`BEQ_rel & T==`Tthree & phi1)
			 | (OP==`BEQ_rel & T==`Tthree & phi2)
			 | (OP==`SBC_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`SBC_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`SBC_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`SBC_izy & T==`TzeroCrossPg & phi2)
			 | (OP==`SBC_izy & T==`Tthree & phi1)
			 | (OP==`SBC_izy & T==`Tthree & phi2)
			 | (OP==`SBC_izy & T==`Tfour & phi1)
			 | (OP==`SBC_izy & T==`Tfour & phi2)
			 | (OP==`SBC_izy & T==`Tfive & phi1)
			 | (OP==`SBC_izy & T==`Tfive & phi2)
			 | (OP==`SBC_zpx & T==`Tzero & phi1)
			 | (OP==`SBC_zpx & T==`Tzero & phi2)
			 | (OP==`SBC_zpx & T==`Tthree & phi1)
			 | (OP==`SBC_zpx & T==`Tthree & phi2)
			 | (OP==`INC_zpx & T==`Tzero & phi1)
			 | (OP==`INC_zpx & T==`Tzero & phi2)
			 | (OP==`INC_zpx & T==`Tthree & phi1)
			 | (OP==`INC_zpx & T==`Tthree & phi2)
			 | (OP==`INC_zpx & T==`Tfour & phi1)
			 | (OP==`INC_zpx & T==`Tfour & phi2)
			 | (OP==`INC_zpx & T==`Tfive & phi1)
			 | (OP==`INC_zpx & T==`Tfive & phi2)
			 | (OP==`SED & T==`Ttwo & phi1)
			 | (OP==`SED & T==`Ttwo & phi2)
			 | (OP==`SBC_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`SBC_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`SBC_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`SBC_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`SBC_aby & T==`Tfour & phi1)
			 | (OP==`SBC_aby & T==`Tfour & phi2)
			 | (OP==`SBC_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`SBC_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`SBC_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`SBC_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`SBC_abx & T==`Tfour & phi1)
			 | (OP==`SBC_abx & T==`Tfour & phi2)
			 | (OP==`INC_abx & T==`Tzero & phi1)
			 | (OP==`INC_abx & T==`Tzero & phi2)
			 | (OP==`INC_abx & T==`Tfour & phi1)
			 | (OP==`INC_abx & T==`Tfour & phi2)
			 | (OP==`INC_abx & T==`Tfive & phi1)
			 | (OP==`INC_abx & T==`Tfive & phi2)
			 | (OP==`INC_abx & T==`Tsix & phi1)
			 | (OP==`INC_abx & T==`Tsix & phi2)
			;

assign control[`PCL_DB] = (OP==`BRK & T==`Tthree & phi2)
			 | (OP==`BRK & T==`Tfour & phi1)
			 | (OP==`JSR_abs & T==`Tfour & phi2)
			 | (OP==`JSR_abs & T==`Tfive & phi1)
			;

assign control[`PCL_ADL] = (OP==`BRK & T==`Tone & phi2)
			 | (OP==`BRK & T==`Ttwo & phi1)
			 | (OP==`ORA_izx & T==`Tzero & phi2)
			 | (OP==`ORA_izx & T==`Tone & phi1)
			 | (OP==`ORA_izx & T==`Tone & phi2)
			 | (OP==`ORA_izx & T==`Ttwo & phi1)
			 | (OP==`ORA_zp & T==`Tzero & phi2)
			 | (OP==`ORA_zp & T==`Tone & phi1)
			 | (OP==`ORA_zp & T==`Tone & phi2)
			 | (OP==`ORA_zp & T==`Ttwo & phi1)
			 | (OP==`ASL_zp & T==`Tzero & phi2)
			 | (OP==`ASL_zp & T==`Tone & phi1)
			 | (OP==`ASL_zp & T==`Tone & phi2)
			 | (OP==`ASL_zp & T==`Ttwo & phi1)
			 | (OP==`PHP & T==`Tzero & phi2)
			 | (OP==`PHP & T==`Tone & phi1)
			 | (OP==`PHP & T==`Tone & phi2)
			 | (OP==`PHP & T==`Ttwo & phi1)
			 | (OP==`ORA_imm & T==`Tone & phi1)
			 | (OP==`ORA_imm & T==`Tone & phi2)
			 | (OP==`ORA_imm & T==`Ttwo & phi1)
			 | (OP==`ORA_imm & T==`Ttwo & phi2)
			 | (OP==`ASL & T==`Tone & phi1)
			 | (OP==`ASL & T==`Tone & phi2)
			 | (OP==`ASL & T==`Ttwo & phi1)
			 | (OP==`ASL & T==`Ttwo & phi2)
			 | (OP==`ORA_abs & T==`Tzero & phi2)
			 | (OP==`ORA_abs & T==`Tone & phi1)
			 | (OP==`ORA_abs & T==`Tone & phi2)
			 | (OP==`ORA_abs & T==`Ttwo & phi1)
			 | (OP==`ORA_abs & T==`Ttwo & phi2)
			 | (OP==`ORA_abs & T==`Tthree & phi1)
			 | (OP==`ASL_abs & T==`Tzero & phi2)
			 | (OP==`ASL_abs & T==`Tone & phi1)
			 | (OP==`ASL_abs & T==`Tone & phi2)
			 | (OP==`ASL_abs & T==`Ttwo & phi1)
			 | (OP==`ASL_abs & T==`Ttwo & phi2)
			 | (OP==`ASL_abs & T==`Tthree & phi1)
			 | (OP==`BPL_rel & T==`Tzero & phi2)
			 | (OP==`BPL_rel & T==`Ttwo & phi1)
			 | (OP==`BPL_rel & T==`Ttwo & phi2)
			 | (OP==`BPL_rel & T==`Tthree & phi1)
			 | (OP==`BPL_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BPL_rel & T==`T1BranchCross & phi1)
			 | (OP==`BPL_rel & T==`T1BranchCross & phi2)
			 | (OP==`BPL_rel & T==`T1NoBranch & phi1)
			 | (OP==`BPL_rel & T==`T1NoBranch & phi2)
			 | (OP==`ORA_izy & T==`TzeroCrossPg & phi2)
			 | (OP==`ORA_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`ORA_izy & T==`Tone & phi1)
			 | (OP==`ORA_izy & T==`Tone & phi2)
			 | (OP==`ORA_izy & T==`Ttwo & phi1)
			 | (OP==`ORA_zpx & T==`Tzero & phi2)
			 | (OP==`ORA_zpx & T==`Tone & phi1)
			 | (OP==`ORA_zpx & T==`Tone & phi2)
			 | (OP==`ORA_zpx & T==`Ttwo & phi1)
			 | (OP==`ASL_zpx & T==`Tzero & phi2)
			 | (OP==`ASL_zpx & T==`Tone & phi1)
			 | (OP==`ASL_zpx & T==`Tone & phi2)
			 | (OP==`ASL_zpx & T==`Ttwo & phi1)
			 | (OP==`CLC & T==`Tone & phi1)
			 | (OP==`CLC & T==`Tone & phi2)
			 | (OP==`CLC & T==`Ttwo & phi1)
			 | (OP==`CLC & T==`Ttwo & phi2)
			 | (OP==`ORA_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`ORA_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`ORA_aby & T==`Tone & phi1)
			 | (OP==`ORA_aby & T==`Tone & phi2)
			 | (OP==`ORA_aby & T==`Ttwo & phi1)
			 | (OP==`ORA_aby & T==`Ttwo & phi2)
			 | (OP==`ORA_aby & T==`Tthree & phi1)
			 | (OP==`ORA_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`ORA_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`ORA_abx & T==`Tone & phi1)
			 | (OP==`ORA_abx & T==`Tone & phi2)
			 | (OP==`ORA_abx & T==`Ttwo & phi1)
			 | (OP==`ORA_abx & T==`Ttwo & phi2)
			 | (OP==`ORA_abx & T==`Tthree & phi1)
			 | (OP==`ASL_abx & T==`Tzero & phi2)
			 | (OP==`ASL_abx & T==`Tone & phi1)
			 | (OP==`ASL_abx & T==`Tone & phi2)
			 | (OP==`ASL_abx & T==`Ttwo & phi1)
			 | (OP==`ASL_abx & T==`Ttwo & phi2)
			 | (OP==`ASL_abx & T==`Tthree & phi1)
			 | (OP==`JSR_abs & T==`Tzero & phi1)
			 | (OP==`JSR_abs & T==`Tone & phi2)
			 | (OP==`JSR_abs & T==`Ttwo & phi1)
			 | (OP==`JSR_abs & T==`Tfive & phi2)
			 | (OP==`AND_izx & T==`Tzero & phi2)
			 | (OP==`AND_izx & T==`Tone & phi1)
			 | (OP==`AND_izx & T==`Tone & phi2)
			 | (OP==`AND_izx & T==`Ttwo & phi1)
			 | (OP==`BIT_zp & T==`Tzero & phi2)
			 | (OP==`BIT_zp & T==`Tone & phi1)
			 | (OP==`BIT_zp & T==`Tone & phi2)
			 | (OP==`BIT_zp & T==`Ttwo & phi1)
			 | (OP==`AND_zp & T==`Tzero & phi2)
			 | (OP==`AND_zp & T==`Tone & phi1)
			 | (OP==`AND_zp & T==`Tone & phi2)
			 | (OP==`AND_zp & T==`Ttwo & phi1)
			 | (OP==`ROL_zp & T==`Tzero & phi2)
			 | (OP==`ROL_zp & T==`Tone & phi1)
			 | (OP==`ROL_zp & T==`Tone & phi2)
			 | (OP==`ROL_zp & T==`Ttwo & phi1)
			 | (OP==`PLP & T==`Tzero & phi2)
			 | (OP==`PLP & T==`Tone & phi1)
			 | (OP==`PLP & T==`Tone & phi2)
			 | (OP==`PLP & T==`Ttwo & phi1)
			 | (OP==`AND_imm & T==`Tone & phi1)
			 | (OP==`AND_imm & T==`Tone & phi2)
			 | (OP==`AND_imm & T==`Ttwo & phi1)
			 | (OP==`AND_imm & T==`Ttwo & phi2)
			 | (OP==`ROL & T==`Tone & phi1)
			 | (OP==`ROL & T==`Tone & phi2)
			 | (OP==`ROL & T==`Ttwo & phi1)
			 | (OP==`ROL & T==`Ttwo & phi2)
			 | (OP==`BIT_abs & T==`Tzero & phi2)
			 | (OP==`BIT_abs & T==`Tone & phi1)
			 | (OP==`BIT_abs & T==`Tone & phi2)
			 | (OP==`BIT_abs & T==`Ttwo & phi1)
			 | (OP==`BIT_abs & T==`Ttwo & phi2)
			 | (OP==`BIT_abs & T==`Tthree & phi1)
			 | (OP==`AND_abs & T==`Tzero & phi2)
			 | (OP==`AND_abs & T==`Tone & phi1)
			 | (OP==`AND_abs & T==`Tone & phi2)
			 | (OP==`AND_abs & T==`Ttwo & phi1)
			 | (OP==`AND_abs & T==`Ttwo & phi2)
			 | (OP==`AND_abs & T==`Tthree & phi1)
			 | (OP==`ROL_abs & T==`Tzero & phi2)
			 | (OP==`ROL_abs & T==`Tone & phi1)
			 | (OP==`ROL_abs & T==`Tone & phi2)
			 | (OP==`ROL_abs & T==`Ttwo & phi1)
			 | (OP==`ROL_abs & T==`Ttwo & phi2)
			 | (OP==`ROL_abs & T==`Tthree & phi1)
			 | (OP==`BMI_rel & T==`Tzero & phi2)
			 | (OP==`BMI_rel & T==`Ttwo & phi1)
			 | (OP==`BMI_rel & T==`Ttwo & phi2)
			 | (OP==`BMI_rel & T==`Tthree & phi1)
			 | (OP==`BMI_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BMI_rel & T==`T1BranchCross & phi1)
			 | (OP==`BMI_rel & T==`T1BranchCross & phi2)
			 | (OP==`BMI_rel & T==`T1NoBranch & phi1)
			 | (OP==`BMI_rel & T==`T1NoBranch & phi2)
			 | (OP==`AND_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`AND_izy & T==`TzeroCrossPg & phi2)
			 | (OP==`AND_izy & T==`Tone & phi1)
			 | (OP==`AND_izy & T==`Tone & phi2)
			 | (OP==`AND_izy & T==`Ttwo & phi1)
			 | (OP==`AND_zpx & T==`Tzero & phi2)
			 | (OP==`AND_zpx & T==`Tone & phi1)
			 | (OP==`AND_zpx & T==`Tone & phi2)
			 | (OP==`AND_zpx & T==`Ttwo & phi1)
			 | (OP==`ROL_zpx & T==`Tzero & phi2)
			 | (OP==`ROL_zpx & T==`Tone & phi1)
			 | (OP==`ROL_zpx & T==`Tone & phi2)
			 | (OP==`ROL_zpx & T==`Ttwo & phi1)
			 | (OP==`SEC & T==`Tone & phi1)
			 | (OP==`SEC & T==`Tone & phi2)
			 | (OP==`SEC & T==`Ttwo & phi1)
			 | (OP==`SEC & T==`Ttwo & phi2)
			 | (OP==`AND_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`AND_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`AND_aby & T==`Tone & phi1)
			 | (OP==`AND_aby & T==`Tone & phi2)
			 | (OP==`AND_aby & T==`Ttwo & phi1)
			 | (OP==`AND_aby & T==`Ttwo & phi2)
			 | (OP==`AND_aby & T==`Tthree & phi1)
			 | (OP==`AND_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`AND_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`AND_abx & T==`Tone & phi1)
			 | (OP==`AND_abx & T==`Tone & phi2)
			 | (OP==`AND_abx & T==`Ttwo & phi1)
			 | (OP==`AND_abx & T==`Ttwo & phi2)
			 | (OP==`AND_abx & T==`Tthree & phi1)
			 | (OP==`ROL_abx & T==`Tzero & phi2)
			 | (OP==`ROL_abx & T==`Tone & phi1)
			 | (OP==`ROL_abx & T==`Tone & phi2)
			 | (OP==`ROL_abx & T==`Ttwo & phi1)
			 | (OP==`ROL_abx & T==`Ttwo & phi2)
			 | (OP==`ROL_abx & T==`Tthree & phi1)
			 | (OP==`RTI & T==`Tone & phi2)
			 | (OP==`RTI & T==`Ttwo & phi1)
			 | (OP==`EOR_izx & T==`Tzero & phi2)
			 | (OP==`EOR_izx & T==`Tone & phi1)
			 | (OP==`EOR_izx & T==`Tone & phi2)
			 | (OP==`EOR_izx & T==`Ttwo & phi1)
			 | (OP==`EOR_zp & T==`Tzero & phi2)
			 | (OP==`EOR_zp & T==`Tone & phi1)
			 | (OP==`EOR_zp & T==`Tone & phi2)
			 | (OP==`EOR_zp & T==`Ttwo & phi1)
			 | (OP==`LSR_zp & T==`Tzero & phi2)
			 | (OP==`LSR_zp & T==`Tone & phi1)
			 | (OP==`LSR_zp & T==`Tone & phi2)
			 | (OP==`LSR_zp & T==`Ttwo & phi1)
			 | (OP==`PHA & T==`Tzero & phi2)
			 | (OP==`PHA & T==`Tone & phi1)
			 | (OP==`PHA & T==`Tone & phi2)
			 | (OP==`PHA & T==`Ttwo & phi1)
			 | (OP==`EOR_imm & T==`Tone & phi1)
			 | (OP==`EOR_imm & T==`Tone & phi2)
			 | (OP==`EOR_imm & T==`Ttwo & phi1)
			 | (OP==`EOR_imm & T==`Ttwo & phi2)
			 | (OP==`LSR & T==`Tone & phi1)
			 | (OP==`LSR & T==`Tone & phi2)
			 | (OP==`LSR & T==`Ttwo & phi1)
			 | (OP==`LSR & T==`Ttwo & phi2)
			 | (OP==`JMP_abs & T==`Tzero & phi1)
			 | (OP==`JMP_abs & T==`Tone & phi2)
			 | (OP==`JMP_abs & T==`Ttwo & phi1)
			 | (OP==`JMP_abs & T==`Ttwo & phi2)
			 | (OP==`EOR_abs & T==`Tzero & phi2)
			 | (OP==`EOR_abs & T==`Tone & phi1)
			 | (OP==`EOR_abs & T==`Tone & phi2)
			 | (OP==`EOR_abs & T==`Ttwo & phi1)
			 | (OP==`EOR_abs & T==`Ttwo & phi2)
			 | (OP==`EOR_abs & T==`Tthree & phi1)
			 | (OP==`LSR_abs & T==`Tzero & phi2)
			 | (OP==`LSR_abs & T==`Tone & phi1)
			 | (OP==`LSR_abs & T==`Tone & phi2)
			 | (OP==`LSR_abs & T==`Ttwo & phi1)
			 | (OP==`LSR_abs & T==`Ttwo & phi2)
			 | (OP==`LSR_abs & T==`Tthree & phi1)
			 | (OP==`BVC_rel & T==`Tzero & phi2)
			 | (OP==`BVC_rel & T==`Ttwo & phi1)
			 | (OP==`BVC_rel & T==`Ttwo & phi2)
			 | (OP==`BVC_rel & T==`Tthree & phi1)
			 | (OP==`BVC_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BVC_rel & T==`T1BranchCross & phi1)
			 | (OP==`BVC_rel & T==`T1BranchCross & phi2)
			 | (OP==`BVC_rel & T==`T1NoBranch & phi1)
			 | (OP==`BVC_rel & T==`T1NoBranch & phi2)
			 | (OP==`EOR_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`EOR_izy & T==`TzeroCrossPg & phi2)
			 | (OP==`EOR_izy & T==`Tone & phi1)
			 | (OP==`EOR_izy & T==`Tone & phi2)
			 | (OP==`EOR_izy & T==`Ttwo & phi1)
			 | (OP==`EOR_zpx & T==`Tzero & phi2)
			 | (OP==`EOR_zpx & T==`Tone & phi1)
			 | (OP==`EOR_zpx & T==`Tone & phi2)
			 | (OP==`EOR_zpx & T==`Ttwo & phi1)
			 | (OP==`LSR_zpx & T==`Tzero & phi2)
			 | (OP==`LSR_zpx & T==`Tone & phi1)
			 | (OP==`LSR_zpx & T==`Tone & phi2)
			 | (OP==`LSR_zpx & T==`Ttwo & phi1)
			 | (OP==`CLI & T==`Tone & phi1)
			 | (OP==`CLI & T==`Tone & phi2)
			 | (OP==`CLI & T==`Ttwo & phi1)
			 | (OP==`CLI & T==`Ttwo & phi2)
			 | (OP==`EOR_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`EOR_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`EOR_aby & T==`Tone & phi1)
			 | (OP==`EOR_aby & T==`Tone & phi2)
			 | (OP==`EOR_aby & T==`Ttwo & phi1)
			 | (OP==`EOR_aby & T==`Ttwo & phi2)
			 | (OP==`EOR_aby & T==`Tthree & phi1)
			 | (OP==`EOR_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`EOR_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`EOR_abx & T==`Tone & phi1)
			 | (OP==`EOR_abx & T==`Tone & phi2)
			 | (OP==`EOR_abx & T==`Ttwo & phi1)
			 | (OP==`EOR_abx & T==`Ttwo & phi2)
			 | (OP==`EOR_abx & T==`Tthree & phi1)
			 | (OP==`LSR_abx & T==`Tzero & phi2)
			 | (OP==`LSR_abx & T==`Tone & phi1)
			 | (OP==`LSR_abx & T==`Tone & phi2)
			 | (OP==`LSR_abx & T==`Ttwo & phi1)
			 | (OP==`LSR_abx & T==`Ttwo & phi2)
			 | (OP==`LSR_abx & T==`Tthree & phi1)
			 | (OP==`RTS & T==`Tzero & phi2)
			 | (OP==`RTS & T==`Tone & phi1)
			 | (OP==`RTS & T==`Tone & phi2)
			 | (OP==`RTS & T==`Ttwo & phi1)
			 | (OP==`ADC_izx & T==`Tzero & phi2)
			 | (OP==`ADC_izx & T==`Tone & phi1)
			 | (OP==`ADC_izx & T==`Tone & phi2)
			 | (OP==`ADC_izx & T==`Ttwo & phi1)
			 | (OP==`ADC_zp & T==`Tzero & phi2)
			 | (OP==`ADC_zp & T==`Tone & phi1)
			 | (OP==`ADC_zp & T==`Tone & phi2)
			 | (OP==`ADC_zp & T==`Ttwo & phi1)
			 | (OP==`ROR_zp & T==`Tzero & phi2)
			 | (OP==`ROR_zp & T==`Tone & phi1)
			 | (OP==`ROR_zp & T==`Tone & phi2)
			 | (OP==`ROR_zp & T==`Ttwo & phi1)
			 | (OP==`PLA & T==`Tzero & phi2)
			 | (OP==`PLA & T==`Tone & phi1)
			 | (OP==`PLA & T==`Tone & phi2)
			 | (OP==`PLA & T==`Ttwo & phi1)
			 | (OP==`ADC_imm & T==`Tone & phi1)
			 | (OP==`ADC_imm & T==`Tone & phi2)
			 | (OP==`ADC_imm & T==`Ttwo & phi1)
			 | (OP==`ADC_imm & T==`Ttwo & phi2)
			 | (OP==`ROR & T==`Tone & phi1)
			 | (OP==`ROR & T==`Tone & phi2)
			 | (OP==`ROR & T==`Ttwo & phi1)
			 | (OP==`ROR & T==`Ttwo & phi2)
			 | (OP==`JMP_zp & T==`Tone & phi2)
			 | (OP==`JMP_zp & T==`Ttwo & phi1)
			 | (OP==`JMP_zp & T==`Ttwo & phi2)
			 | (OP==`JMP_zp & T==`Tthree & phi1)
			 | (OP==`ADC_abs & T==`Tzero & phi2)
			 | (OP==`ADC_abs & T==`Tone & phi1)
			 | (OP==`ADC_abs & T==`Tone & phi2)
			 | (OP==`ADC_abs & T==`Ttwo & phi1)
			 | (OP==`ADC_abs & T==`Ttwo & phi2)
			 | (OP==`ADC_abs & T==`Tthree & phi1)
			 | (OP==`ROR_abs & T==`Tzero & phi2)
			 | (OP==`ROR_abs & T==`Tone & phi1)
			 | (OP==`ROR_abs & T==`Tone & phi2)
			 | (OP==`ROR_abs & T==`Ttwo & phi1)
			 | (OP==`ROR_abs & T==`Ttwo & phi2)
			 | (OP==`ROR_abs & T==`Tthree & phi1)
			 | (OP==`BVS_rel & T==`Tzero & phi2)
			 | (OP==`BVS_rel & T==`Ttwo & phi1)
			 | (OP==`BVS_rel & T==`Ttwo & phi2)
			 | (OP==`BVS_rel & T==`Tthree & phi1)
			 | (OP==`BVS_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BVS_rel & T==`T1BranchCross & phi1)
			 | (OP==`BVS_rel & T==`T1BranchCross & phi2)
			 | (OP==`BVS_rel & T==`T1NoBranch & phi1)
			 | (OP==`BVS_rel & T==`T1NoBranch & phi2)
			 | (OP==`ADC_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`ADC_izy & T==`TzeroCrossPg & phi2)
			 | (OP==`ADC_izy & T==`Tone & phi1)
			 | (OP==`ADC_izy & T==`Tone & phi2)
			 | (OP==`ADC_izy & T==`Ttwo & phi1)
			 | (OP==`ADC_zpx & T==`Tzero & phi2)
			 | (OP==`ADC_zpx & T==`Tone & phi1)
			 | (OP==`ADC_zpx & T==`Tone & phi2)
			 | (OP==`ADC_zpx & T==`Ttwo & phi1)
			 | (OP==`ROR_zpx & T==`Tzero & phi2)
			 | (OP==`ROR_zpx & T==`Tone & phi1)
			 | (OP==`ROR_zpx & T==`Tone & phi2)
			 | (OP==`ROR_zpx & T==`Ttwo & phi1)
			 | (OP==`SEI & T==`Tone & phi1)
			 | (OP==`SEI & T==`Tone & phi2)
			 | (OP==`SEI & T==`Ttwo & phi1)
			 | (OP==`SEI & T==`Ttwo & phi2)
			 | (OP==`ADC_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`ADC_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`ADC_aby & T==`Tone & phi1)
			 | (OP==`ADC_aby & T==`Tone & phi2)
			 | (OP==`ADC_aby & T==`Ttwo & phi1)
			 | (OP==`ADC_aby & T==`Ttwo & phi2)
			 | (OP==`ADC_aby & T==`Tthree & phi1)
			 | (OP==`ADC_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`ADC_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`ADC_abx & T==`Tone & phi1)
			 | (OP==`ADC_abx & T==`Tone & phi2)
			 | (OP==`ADC_abx & T==`Ttwo & phi1)
			 | (OP==`ADC_abx & T==`Ttwo & phi2)
			 | (OP==`ADC_abx & T==`Tthree & phi1)
			 | (OP==`ROR_abx & T==`Tzero & phi2)
			 | (OP==`ROR_abx & T==`Tone & phi1)
			 | (OP==`ROR_abx & T==`Tone & phi2)
			 | (OP==`ROR_abx & T==`Ttwo & phi1)
			 | (OP==`ROR_abx & T==`Ttwo & phi2)
			 | (OP==`ROR_abx & T==`Tthree & phi1)
			 | (OP==`STA_izx & T==`Tzero & phi2)
			 | (OP==`STA_izx & T==`Tone & phi1)
			 | (OP==`STA_izx & T==`Tone & phi2)
			 | (OP==`STA_izx & T==`Ttwo & phi1)
			 | (OP==`STY_zp & T==`Tzero & phi2)
			 | (OP==`STY_zp & T==`Tone & phi1)
			 | (OP==`STY_zp & T==`Tone & phi2)
			 | (OP==`STY_zp & T==`Ttwo & phi1)
			 | (OP==`STA_zp & T==`Tzero & phi2)
			 | (OP==`STA_zp & T==`Tone & phi1)
			 | (OP==`STA_zp & T==`Tone & phi2)
			 | (OP==`STA_zp & T==`Ttwo & phi1)
			 | (OP==`STX_zp & T==`Tzero & phi2)
			 | (OP==`STX_zp & T==`Tone & phi1)
			 | (OP==`STX_zp & T==`Tone & phi2)
			 | (OP==`STX_zp & T==`Ttwo & phi1)
			 | (OP==`DEY & T==`Tone & phi1)
			 | (OP==`DEY & T==`Tone & phi2)
			 | (OP==`DEY & T==`Ttwo & phi1)
			 | (OP==`DEY & T==`Ttwo & phi2)
			 | (OP==`TXA & T==`Tone & phi1)
			 | (OP==`TXA & T==`Tone & phi2)
			 | (OP==`TXA & T==`Ttwo & phi1)
			 | (OP==`TXA & T==`Ttwo & phi2)
			 | (OP==`STY_abs & T==`Tzero & phi2)
			 | (OP==`STY_abs & T==`Tone & phi1)
			 | (OP==`STY_abs & T==`Tone & phi2)
			 | (OP==`STY_abs & T==`Ttwo & phi1)
			 | (OP==`STY_abs & T==`Ttwo & phi2)
			 | (OP==`STY_abs & T==`Tthree & phi1)
			 | (OP==`STA_abs & T==`Tzero & phi2)
			 | (OP==`STA_abs & T==`Tone & phi1)
			 | (OP==`STA_abs & T==`Tone & phi2)
			 | (OP==`STA_abs & T==`Ttwo & phi1)
			 | (OP==`STA_abs & T==`Ttwo & phi2)
			 | (OP==`STA_abs & T==`Tthree & phi1)
			 | (OP==`STX_abs & T==`Tzero & phi2)
			 | (OP==`STX_abs & T==`Tone & phi1)
			 | (OP==`STX_abs & T==`Tone & phi2)
			 | (OP==`STX_abs & T==`Ttwo & phi1)
			 | (OP==`STX_abs & T==`Ttwo & phi2)
			 | (OP==`STX_abs & T==`Tthree & phi1)
			 | (OP==`BCC_rel & T==`Tzero & phi2)
			 | (OP==`BCC_rel & T==`Ttwo & phi1)
			 | (OP==`BCC_rel & T==`Ttwo & phi2)
			 | (OP==`BCC_rel & T==`Tthree & phi1)
			 | (OP==`BCC_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BCC_rel & T==`T1BranchCross & phi1)
			 | (OP==`BCC_rel & T==`T1BranchCross & phi2)
			 | (OP==`BCC_rel & T==`T1NoBranch & phi1)
			 | (OP==`BCC_rel & T==`T1NoBranch & phi2)
			 | (OP==`STA_izy & T==`Tzero & phi2)
			 | (OP==`STA_izy & T==`Tone & phi1)
			 | (OP==`STA_izy & T==`Tone & phi2)
			 | (OP==`STA_izy & T==`Ttwo & phi1)
			 | (OP==`STY_zpx & T==`Tzero & phi2)
			 | (OP==`STY_zpx & T==`Tone & phi1)
			 | (OP==`STY_zpx & T==`Tone & phi2)
			 | (OP==`STY_zpx & T==`Ttwo & phi1)
			 | (OP==`STA_zpx & T==`Tzero & phi2)
			 | (OP==`STA_zpx & T==`Tone & phi1)
			 | (OP==`STA_zpx & T==`Tone & phi2)
			 | (OP==`STA_zpx & T==`Ttwo & phi1)
			 | (OP==`STX_zpy & T==`Tzero & phi2)
			 | (OP==`STX_zpy & T==`Tone & phi1)
			 | (OP==`STX_zpy & T==`Tone & phi2)
			 | (OP==`STX_zpy & T==`Ttwo & phi1)
			 | (OP==`TYA & T==`Tone & phi1)
			 | (OP==`TYA & T==`Tone & phi2)
			 | (OP==`TYA & T==`Ttwo & phi1)
			 | (OP==`TYA & T==`Ttwo & phi2)
			 | (OP==`STA_aby & T==`Tzero & phi2)
			 | (OP==`STA_aby & T==`Tone & phi1)
			 | (OP==`STA_aby & T==`Tone & phi2)
			 | (OP==`STA_aby & T==`Ttwo & phi1)
			 | (OP==`STA_aby & T==`Ttwo & phi2)
			 | (OP==`STA_aby & T==`Tthree & phi1)
			 | (OP==`TXS & T==`Tone & phi1)
			 | (OP==`TXS & T==`Tone & phi2)
			 | (OP==`TXS & T==`Ttwo & phi1)
			 | (OP==`TXS & T==`Ttwo & phi2)
			 | (OP==`STA_abx & T==`Tzero & phi2)
			 | (OP==`STA_abx & T==`Tone & phi1)
			 | (OP==`STA_abx & T==`Tone & phi2)
			 | (OP==`STA_abx & T==`Ttwo & phi1)
			 | (OP==`STA_abx & T==`Ttwo & phi2)
			 | (OP==`STA_abx & T==`Tthree & phi1)
			 | (OP==`LDY_imm & T==`Tone & phi1)
			 | (OP==`LDY_imm & T==`Tone & phi2)
			 | (OP==`LDY_imm & T==`Ttwo & phi1)
			 | (OP==`LDY_imm & T==`Ttwo & phi2)
			 | (OP==`LDA_izx & T==`Tzero & phi2)
			 | (OP==`LDA_izx & T==`Tone & phi1)
			 | (OP==`LDA_izx & T==`Tone & phi2)
			 | (OP==`LDA_izx & T==`Ttwo & phi1)
			 | (OP==`LDX_imm & T==`Tone & phi1)
			 | (OP==`LDX_imm & T==`Tone & phi2)
			 | (OP==`LDX_imm & T==`Ttwo & phi1)
			 | (OP==`LDX_imm & T==`Ttwo & phi2)
			 | (OP==`LDY_zp & T==`Tzero & phi2)
			 | (OP==`LDY_zp & T==`Tone & phi1)
			 | (OP==`LDY_zp & T==`Tone & phi2)
			 | (OP==`LDY_zp & T==`Ttwo & phi1)
			 | (OP==`LDA_zp & T==`Tzero & phi2)
			 | (OP==`LDA_zp & T==`Tone & phi1)
			 | (OP==`LDA_zp & T==`Tone & phi2)
			 | (OP==`LDA_zp & T==`Ttwo & phi1)
			 | (OP==`LDX_zp & T==`Tzero & phi2)
			 | (OP==`LDX_zp & T==`Tone & phi1)
			 | (OP==`LDX_zp & T==`Tone & phi2)
			 | (OP==`LDX_zp & T==`Ttwo & phi1)
			 | (OP==`TAY & T==`Tone & phi1)
			 | (OP==`TAY & T==`Tone & phi2)
			 | (OP==`TAY & T==`Ttwo & phi1)
			 | (OP==`TAY & T==`Ttwo & phi2)
			 | (OP==`LDA_imm & T==`Tone & phi1)
			 | (OP==`LDA_imm & T==`Tone & phi2)
			 | (OP==`LDA_imm & T==`Ttwo & phi1)
			 | (OP==`LDA_imm & T==`Ttwo & phi2)
			 | (OP==`TAX & T==`Tone & phi1)
			 | (OP==`TAX & T==`Tone & phi2)
			 | (OP==`TAX & T==`Ttwo & phi1)
			 | (OP==`TAX & T==`Ttwo & phi2)
			 | (OP==`LDY_abs & T==`Tzero & phi2)
			 | (OP==`LDY_abs & T==`Tone & phi1)
			 | (OP==`LDY_abs & T==`Tone & phi2)
			 | (OP==`LDY_abs & T==`Ttwo & phi1)
			 | (OP==`LDY_abs & T==`Ttwo & phi2)
			 | (OP==`LDY_abs & T==`Tthree & phi1)
			 | (OP==`LDA_abs & T==`Tzero & phi2)
			 | (OP==`LDA_abs & T==`Tone & phi1)
			 | (OP==`LDA_abs & T==`Tone & phi2)
			 | (OP==`LDA_abs & T==`Ttwo & phi1)
			 | (OP==`LDA_abs & T==`Ttwo & phi2)
			 | (OP==`LDA_abs & T==`Tthree & phi1)
			 | (OP==`LDX_abs & T==`Tzero & phi2)
			 | (OP==`LDX_abs & T==`Tone & phi1)
			 | (OP==`LDX_abs & T==`Tone & phi2)
			 | (OP==`LDX_abs & T==`Ttwo & phi1)
			 | (OP==`LDX_abs & T==`Ttwo & phi2)
			 | (OP==`LDX_abs & T==`Tthree & phi1)
			 | (OP==`BCS_rel & T==`Tzero & phi2)
			 | (OP==`BCS_rel & T==`Ttwo & phi1)
			 | (OP==`BCS_rel & T==`Ttwo & phi2)
			 | (OP==`BCS_rel & T==`Tthree & phi1)
			 | (OP==`BCS_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BCS_rel & T==`T1BranchCross & phi1)
			 | (OP==`BCS_rel & T==`T1BranchCross & phi2)
			 | (OP==`BCS_rel & T==`T1NoBranch & phi1)
			 | (OP==`BCS_rel & T==`T1NoBranch & phi2)
			 | (OP==`LDA_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`LDA_izy & T==`TzeroCrossPg & phi2)
			 | (OP==`LDA_izy & T==`Tone & phi1)
			 | (OP==`LDA_izy & T==`Tone & phi2)
			 | (OP==`LDA_izy & T==`Ttwo & phi1)
			 | (OP==`LDY_zpx & T==`Tzero & phi2)
			 | (OP==`LDY_zpx & T==`Tone & phi1)
			 | (OP==`LDY_zpx & T==`Tone & phi2)
			 | (OP==`LDY_zpx & T==`Ttwo & phi1)
			 | (OP==`LDA_zpx & T==`Tzero & phi2)
			 | (OP==`LDA_zpx & T==`Tone & phi1)
			 | (OP==`LDA_zpx & T==`Tone & phi2)
			 | (OP==`LDA_zpx & T==`Ttwo & phi1)
			 | (OP==`LDX_zpy & T==`Tzero & phi2)
			 | (OP==`LDX_zpy & T==`Tone & phi1)
			 | (OP==`LDX_zpy & T==`Tone & phi2)
			 | (OP==`LDX_zpy & T==`Ttwo & phi1)
			 | (OP==`CLV & T==`Tone & phi1)
			 | (OP==`CLV & T==`Tone & phi2)
			 | (OP==`CLV & T==`Ttwo & phi1)
			 | (OP==`CLV & T==`Ttwo & phi2)
			 | (OP==`LDA_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`LDA_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`LDA_aby & T==`Tone & phi1)
			 | (OP==`LDA_aby & T==`Tone & phi2)
			 | (OP==`LDA_aby & T==`Ttwo & phi1)
			 | (OP==`LDA_aby & T==`Ttwo & phi2)
			 | (OP==`LDA_aby & T==`Tthree & phi1)
			 | (OP==`TSX & T==`Tone & phi1)
			 | (OP==`TSX & T==`Tone & phi2)
			 | (OP==`TSX & T==`Ttwo & phi1)
			 | (OP==`TSX & T==`Ttwo & phi2)
			 | (OP==`LDY_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`LDY_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`LDY_abx & T==`Tone & phi1)
			 | (OP==`LDY_abx & T==`Tone & phi2)
			 | (OP==`LDY_abx & T==`Ttwo & phi1)
			 | (OP==`LDY_abx & T==`Ttwo & phi2)
			 | (OP==`LDY_abx & T==`Tthree & phi1)
			 | (OP==`LDA_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`LDA_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`LDA_abx & T==`Tone & phi1)
			 | (OP==`LDA_abx & T==`Tone & phi2)
			 | (OP==`LDA_abx & T==`Ttwo & phi1)
			 | (OP==`LDA_abx & T==`Ttwo & phi2)
			 | (OP==`LDA_abx & T==`Tthree & phi1)
			 | (OP==`LDX_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`LDX_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`LDX_aby & T==`Tone & phi1)
			 | (OP==`LDX_aby & T==`Tone & phi2)
			 | (OP==`LDX_aby & T==`Ttwo & phi1)
			 | (OP==`LDX_aby & T==`Ttwo & phi2)
			 | (OP==`LDX_aby & T==`Tthree & phi1)
			 | (OP==`CPY_imm & T==`Tone & phi1)
			 | (OP==`CPY_imm & T==`Tone & phi2)
			 | (OP==`CPY_imm & T==`Ttwo & phi1)
			 | (OP==`CPY_imm & T==`Ttwo & phi2)
			 | (OP==`CMP_izx & T==`Tzero & phi2)
			 | (OP==`CMP_izx & T==`Tone & phi1)
			 | (OP==`CMP_izx & T==`Tone & phi2)
			 | (OP==`CMP_izx & T==`Ttwo & phi1)
			 | (OP==`CPY_zp & T==`Tzero & phi2)
			 | (OP==`CPY_zp & T==`Tone & phi1)
			 | (OP==`CPY_zp & T==`Tone & phi2)
			 | (OP==`CPY_zp & T==`Ttwo & phi1)
			 | (OP==`CMP_zp & T==`Tzero & phi2)
			 | (OP==`CMP_zp & T==`Tone & phi1)
			 | (OP==`CMP_zp & T==`Tone & phi2)
			 | (OP==`CMP_zp & T==`Ttwo & phi1)
			 | (OP==`DEC_zp & T==`Tzero & phi2)
			 | (OP==`DEC_zp & T==`Tone & phi1)
			 | (OP==`DEC_zp & T==`Tone & phi2)
			 | (OP==`DEC_zp & T==`Ttwo & phi1)
			 | (OP==`INY & T==`Tone & phi1)
			 | (OP==`INY & T==`Tone & phi2)
			 | (OP==`INY & T==`Ttwo & phi1)
			 | (OP==`INY & T==`Ttwo & phi2)
			 | (OP==`CMP_imm & T==`Tone & phi1)
			 | (OP==`CMP_imm & T==`Tone & phi2)
			 | (OP==`CMP_imm & T==`Ttwo & phi1)
			 | (OP==`CMP_imm & T==`Ttwo & phi2)
			 | (OP==`DEX & T==`Tone & phi1)
			 | (OP==`DEX & T==`Tone & phi2)
			 | (OP==`DEX & T==`Ttwo & phi1)
			 | (OP==`DEX & T==`Ttwo & phi2)
			 | (OP==`CPY_abs & T==`Tzero & phi2)
			 | (OP==`CPY_abs & T==`Tone & phi1)
			 | (OP==`CPY_abs & T==`Tone & phi2)
			 | (OP==`CPY_abs & T==`Ttwo & phi1)
			 | (OP==`CPY_abs & T==`Ttwo & phi2)
			 | (OP==`CPY_abs & T==`Tthree & phi1)
			 | (OP==`CMP_abs & T==`Tzero & phi2)
			 | (OP==`CMP_abs & T==`Tone & phi1)
			 | (OP==`CMP_abs & T==`Tone & phi2)
			 | (OP==`CMP_abs & T==`Ttwo & phi1)
			 | (OP==`CMP_abs & T==`Ttwo & phi2)
			 | (OP==`CMP_abs & T==`Tthree & phi1)
			 | (OP==`DEC_abs & T==`Tzero & phi2)
			 | (OP==`DEC_abs & T==`Tone & phi1)
			 | (OP==`DEC_abs & T==`Tone & phi2)
			 | (OP==`DEC_abs & T==`Ttwo & phi1)
			 | (OP==`DEC_abs & T==`Ttwo & phi2)
			 | (OP==`DEC_abs & T==`Tthree & phi1)
			 | (OP==`BNE_rel & T==`Tzero & phi2)
			 | (OP==`BNE_rel & T==`Ttwo & phi1)
			 | (OP==`BNE_rel & T==`Ttwo & phi2)
			 | (OP==`BNE_rel & T==`Tthree & phi1)
			 | (OP==`BNE_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BNE_rel & T==`T1BranchCross & phi1)
			 | (OP==`BNE_rel & T==`T1BranchCross & phi2)
			 | (OP==`BNE_rel & T==`T1NoBranch & phi1)
			 | (OP==`BNE_rel & T==`T1NoBranch & phi2)
			 | (OP==`CMP_izy & T==`TzeroCrossPg & phi2)
			 | (OP==`CMP_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`CMP_izy & T==`Tone & phi1)
			 | (OP==`CMP_izy & T==`Tone & phi2)
			 | (OP==`CMP_izy & T==`Ttwo & phi1)
			 | (OP==`CMP_zpx & T==`Tzero & phi2)
			 | (OP==`CMP_zpx & T==`Tone & phi1)
			 | (OP==`CMP_zpx & T==`Tone & phi2)
			 | (OP==`CMP_zpx & T==`Ttwo & phi1)
			 | (OP==`DEC_zpx & T==`Tzero & phi2)
			 | (OP==`DEC_zpx & T==`Tone & phi1)
			 | (OP==`DEC_zpx & T==`Tone & phi2)
			 | (OP==`DEC_zpx & T==`Ttwo & phi1)
			 | (OP==`CLD & T==`Tone & phi1)
			 | (OP==`CLD & T==`Tone & phi2)
			 | (OP==`CLD & T==`Ttwo & phi1)
			 | (OP==`CLD & T==`Ttwo & phi2)
			 | (OP==`CMP_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`CMP_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`CMP_aby & T==`Tone & phi1)
			 | (OP==`CMP_aby & T==`Tone & phi2)
			 | (OP==`CMP_aby & T==`Ttwo & phi1)
			 | (OP==`CMP_aby & T==`Ttwo & phi2)
			 | (OP==`CMP_aby & T==`Tthree & phi1)
			 | (OP==`CMP_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`CMP_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`CMP_abx & T==`Tone & phi1)
			 | (OP==`CMP_abx & T==`Tone & phi2)
			 | (OP==`CMP_abx & T==`Ttwo & phi1)
			 | (OP==`CMP_abx & T==`Ttwo & phi2)
			 | (OP==`CMP_abx & T==`Tthree & phi1)
			 | (OP==`DEC_abx & T==`Tzero & phi2)
			 | (OP==`DEC_abx & T==`Tone & phi1)
			 | (OP==`DEC_abx & T==`Tone & phi2)
			 | (OP==`DEC_abx & T==`Ttwo & phi1)
			 | (OP==`DEC_abx & T==`Ttwo & phi2)
			 | (OP==`DEC_abx & T==`Tthree & phi1)
			 | (OP==`CPX_imm & T==`Tone & phi1)
			 | (OP==`CPX_imm & T==`Tone & phi2)
			 | (OP==`CPX_imm & T==`Ttwo & phi1)
			 | (OP==`CPX_imm & T==`Ttwo & phi2)
			 | (OP==`SBC_izx & T==`Tzero & phi2)
			 | (OP==`SBC_izx & T==`Tone & phi1)
			 | (OP==`SBC_izx & T==`Tone & phi2)
			 | (OP==`SBC_izx & T==`Ttwo & phi1)
			 | (OP==`CPX_zp & T==`Tzero & phi2)
			 | (OP==`CPX_zp & T==`Tone & phi1)
			 | (OP==`CPX_zp & T==`Tone & phi2)
			 | (OP==`CPX_zp & T==`Ttwo & phi1)
			 | (OP==`SBC_zp & T==`Tzero & phi2)
			 | (OP==`SBC_zp & T==`Tone & phi1)
			 | (OP==`SBC_zp & T==`Tone & phi2)
			 | (OP==`SBC_zp & T==`Ttwo & phi1)
			 | (OP==`INC_zp & T==`Tzero & phi2)
			 | (OP==`INC_zp & T==`Tone & phi1)
			 | (OP==`INC_zp & T==`Tone & phi2)
			 | (OP==`INC_zp & T==`Ttwo & phi1)
			 | (OP==`INX & T==`Tone & phi1)
			 | (OP==`INX & T==`Tone & phi2)
			 | (OP==`INX & T==`Ttwo & phi1)
			 | (OP==`INX & T==`Ttwo & phi2)
			 | (OP==`SBC_imm & T==`Tone & phi1)
			 | (OP==`SBC_imm & T==`Tone & phi2)
			 | (OP==`SBC_imm & T==`Ttwo & phi1)
			 | (OP==`SBC_imm & T==`Ttwo & phi2)
			 | (OP==`NOP & T==`Tone & phi1)
			 | (OP==`NOP & T==`Tone & phi2)
			 | (OP==`NOP & T==`Ttwo & phi1)
			 | (OP==`NOP & T==`Ttwo & phi2)
			 | (OP==`CPX_abs & T==`Tzero & phi2)
			 | (OP==`CPX_abs & T==`Tone & phi1)
			 | (OP==`CPX_abs & T==`Tone & phi2)
			 | (OP==`CPX_abs & T==`Ttwo & phi1)
			 | (OP==`CPX_abs & T==`Ttwo & phi2)
			 | (OP==`CPX_abs & T==`Tthree & phi1)
			 | (OP==`SBC_abs & T==`Tzero & phi2)
			 | (OP==`SBC_abs & T==`Tone & phi1)
			 | (OP==`SBC_abs & T==`Tone & phi2)
			 | (OP==`SBC_abs & T==`Ttwo & phi1)
			 | (OP==`SBC_abs & T==`Ttwo & phi2)
			 | (OP==`SBC_abs & T==`Tthree & phi1)
			 | (OP==`INC_abs & T==`Tzero & phi2)
			 | (OP==`INC_abs & T==`Tone & phi1)
			 | (OP==`INC_abs & T==`Tone & phi2)
			 | (OP==`INC_abs & T==`Ttwo & phi1)
			 | (OP==`INC_abs & T==`Ttwo & phi2)
			 | (OP==`INC_abs & T==`Tthree & phi1)
			 | (OP==`BEQ_rel & T==`Tzero & phi2)
			 | (OP==`BEQ_rel & T==`Ttwo & phi1)
			 | (OP==`BEQ_rel & T==`Ttwo & phi2)
			 | (OP==`BEQ_rel & T==`Tthree & phi1)
			 | (OP==`BEQ_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BEQ_rel & T==`T1BranchCross & phi1)
			 | (OP==`BEQ_rel & T==`T1BranchCross & phi2)
			 | (OP==`BEQ_rel & T==`T1NoBranch & phi1)
			 | (OP==`BEQ_rel & T==`T1NoBranch & phi2)
			 | (OP==`SBC_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`SBC_izy & T==`TzeroCrossPg & phi2)
			 | (OP==`SBC_izy & T==`Tone & phi1)
			 | (OP==`SBC_izy & T==`Tone & phi2)
			 | (OP==`SBC_izy & T==`Ttwo & phi1)
			 | (OP==`SBC_zpx & T==`Tzero & phi2)
			 | (OP==`SBC_zpx & T==`Tone & phi1)
			 | (OP==`SBC_zpx & T==`Tone & phi2)
			 | (OP==`SBC_zpx & T==`Ttwo & phi1)
			 | (OP==`INC_zpx & T==`Tzero & phi2)
			 | (OP==`INC_zpx & T==`Tone & phi1)
			 | (OP==`INC_zpx & T==`Tone & phi2)
			 | (OP==`INC_zpx & T==`Ttwo & phi1)
			 | (OP==`SED & T==`Tone & phi1)
			 | (OP==`SED & T==`Tone & phi2)
			 | (OP==`SED & T==`Ttwo & phi1)
			 | (OP==`SED & T==`Ttwo & phi2)
			 | (OP==`SBC_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`SBC_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`SBC_aby & T==`Tone & phi1)
			 | (OP==`SBC_aby & T==`Tone & phi2)
			 | (OP==`SBC_aby & T==`Ttwo & phi1)
			 | (OP==`SBC_aby & T==`Ttwo & phi2)
			 | (OP==`SBC_aby & T==`Tthree & phi1)
			 | (OP==`SBC_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`SBC_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`SBC_abx & T==`Tone & phi1)
			 | (OP==`SBC_abx & T==`Tone & phi2)
			 | (OP==`SBC_abx & T==`Ttwo & phi1)
			 | (OP==`SBC_abx & T==`Ttwo & phi2)
			 | (OP==`SBC_abx & T==`Tthree & phi1)
			 | (OP==`INC_abx & T==`Tzero & phi2)
			 | (OP==`INC_abx & T==`Tone & phi1)
			 | (OP==`INC_abx & T==`Tone & phi2)
			 | (OP==`INC_abx & T==`Ttwo & phi1)
			 | (OP==`INC_abx & T==`Ttwo & phi2)
			 | (OP==`INC_abx & T==`Tthree & phi1)
			;

assign control[`PCH_PCH] = (OP==`BRK & T==`Tzero & phi1)
			 | (OP==`BRK & T==`Tthree & phi1)
			 | (OP==`BRK & T==`Tfour & phi1)
			 | (OP==`BRK & T==`Tfive & phi1)
			 | (OP==`BRK & T==`Tsix & phi1)
			 | (OP==`ORA_izx & T==`Tzero & phi1)
			 | (OP==`ORA_izx & T==`Tthree & phi1)
			 | (OP==`ORA_izx & T==`Tfour & phi1)
			 | (OP==`ORA_izx & T==`Tfive & phi1)
			 | (OP==`ORA_zp & T==`Tzero & phi1)
			 | (OP==`ASL_zp & T==`Tzero & phi1)
			 | (OP==`ASL_zp & T==`Tthree & phi1)
			 | (OP==`ASL_zp & T==`Tfour & phi1)
			 | (OP==`PHP & T==`Tzero & phi1)
			 | (OP==`ORA_abs & T==`Tzero & phi1)
			 | (OP==`ASL_abs & T==`Tzero & phi1)
			 | (OP==`ASL_abs & T==`Tfour & phi1)
			 | (OP==`ASL_abs & T==`Tfive & phi1)
			 | (OP==`ORA_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`ORA_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ORA_izy & T==`Tthree & phi1)
			 | (OP==`ORA_izy & T==`Tfour & phi1)
			 | (OP==`ORA_izy & T==`Tfive & phi1)
			 | (OP==`ORA_zpx & T==`Tzero & phi1)
			 | (OP==`ORA_zpx & T==`Tthree & phi1)
			 | (OP==`ASL_zpx & T==`Tzero & phi1)
			 | (OP==`ASL_zpx & T==`Tthree & phi1)
			 | (OP==`ASL_zpx & T==`Tfour & phi1)
			 | (OP==`ASL_zpx & T==`Tfive & phi1)
			 | (OP==`ORA_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ORA_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`ORA_aby & T==`Tfour & phi1)
			 | (OP==`ORA_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ORA_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`ORA_abx & T==`Tfour & phi1)
			 | (OP==`ASL_abx & T==`Tzero & phi1)
			 | (OP==`ASL_abx & T==`Tfour & phi1)
			 | (OP==`ASL_abx & T==`Tfive & phi1)
			 | (OP==`ASL_abx & T==`Tsix & phi1)
			 | (OP==`JSR_abs & T==`Tzero & phi1)
			 | (OP==`JSR_abs & T==`Tthree & phi1)
			 | (OP==`JSR_abs & T==`Tfour & phi1)
			 | (OP==`JSR_abs & T==`Tfive & phi1)
			 | (OP==`AND_izx & T==`Tzero & phi1)
			 | (OP==`AND_izx & T==`Tthree & phi1)
			 | (OP==`AND_izx & T==`Tfour & phi1)
			 | (OP==`AND_izx & T==`Tfive & phi1)
			 | (OP==`BIT_zp & T==`Tzero & phi1)
			 | (OP==`AND_zp & T==`Tzero & phi1)
			 | (OP==`ROL_zp & T==`Tzero & phi1)
			 | (OP==`ROL_zp & T==`Tthree & phi1)
			 | (OP==`ROL_zp & T==`Tfour & phi1)
			 | (OP==`PLP & T==`Tzero & phi1)
			 | (OP==`PLP & T==`Tthree & phi1)
			 | (OP==`BIT_abs & T==`Tzero & phi1)
			 | (OP==`AND_abs & T==`Tzero & phi1)
			 | (OP==`ROL_abs & T==`Tzero & phi1)
			 | (OP==`ROL_abs & T==`Tfour & phi1)
			 | (OP==`ROL_abs & T==`Tfive & phi1)
			 | (OP==`AND_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`AND_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`AND_izy & T==`Tthree & phi1)
			 | (OP==`AND_izy & T==`Tfour & phi1)
			 | (OP==`AND_izy & T==`Tfive & phi1)
			 | (OP==`AND_zpx & T==`Tzero & phi1)
			 | (OP==`AND_zpx & T==`Tthree & phi1)
			 | (OP==`ROL_zpx & T==`Tzero & phi1)
			 | (OP==`ROL_zpx & T==`Tthree & phi1)
			 | (OP==`ROL_zpx & T==`Tfour & phi1)
			 | (OP==`ROL_zpx & T==`Tfive & phi1)
			 | (OP==`AND_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`AND_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`AND_aby & T==`Tfour & phi1)
			 | (OP==`AND_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`AND_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`AND_abx & T==`Tfour & phi1)
			 | (OP==`ROL_abx & T==`Tzero & phi1)
			 | (OP==`ROL_abx & T==`Tfour & phi1)
			 | (OP==`ROL_abx & T==`Tfive & phi1)
			 | (OP==`ROL_abx & T==`Tsix & phi1)
			 | (OP==`RTI & T==`Tzero & phi1)
			 | (OP==`RTI & T==`Tthree & phi1)
			 | (OP==`RTI & T==`Tfour & phi1)
			 | (OP==`RTI & T==`Tfive & phi1)
			 | (OP==`EOR_izx & T==`Tzero & phi1)
			 | (OP==`EOR_izx & T==`Tthree & phi1)
			 | (OP==`EOR_izx & T==`Tfour & phi1)
			 | (OP==`EOR_izx & T==`Tfive & phi1)
			 | (OP==`EOR_zp & T==`Tzero & phi1)
			 | (OP==`LSR_zp & T==`Tzero & phi1)
			 | (OP==`LSR_zp & T==`Tthree & phi1)
			 | (OP==`LSR_zp & T==`Tfour & phi1)
			 | (OP==`PHA & T==`Tzero & phi1)
			 | (OP==`EOR_abs & T==`Tzero & phi1)
			 | (OP==`LSR_abs & T==`Tzero & phi1)
			 | (OP==`LSR_abs & T==`Tfour & phi1)
			 | (OP==`LSR_abs & T==`Tfive & phi1)
			 | (OP==`EOR_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`EOR_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`EOR_izy & T==`Tthree & phi1)
			 | (OP==`EOR_izy & T==`Tfour & phi1)
			 | (OP==`EOR_izy & T==`Tfive & phi1)
			 | (OP==`EOR_zpx & T==`Tzero & phi1)
			 | (OP==`EOR_zpx & T==`Tthree & phi1)
			 | (OP==`LSR_zpx & T==`Tzero & phi1)
			 | (OP==`LSR_zpx & T==`Tthree & phi1)
			 | (OP==`LSR_zpx & T==`Tfour & phi1)
			 | (OP==`LSR_zpx & T==`Tfive & phi1)
			 | (OP==`EOR_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`EOR_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`EOR_aby & T==`Tfour & phi1)
			 | (OP==`EOR_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`EOR_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`EOR_abx & T==`Tfour & phi1)
			 | (OP==`LSR_abx & T==`Tzero & phi1)
			 | (OP==`LSR_abx & T==`Tfour & phi1)
			 | (OP==`LSR_abx & T==`Tfive & phi1)
			 | (OP==`LSR_abx & T==`Tsix & phi1)
			 | (OP==`RTS & T==`Tthree & phi1)
			 | (OP==`RTS & T==`Tfour & phi1)
			 | (OP==`RTS & T==`Tfive & phi1)
			 | (OP==`ADC_izx & T==`Tzero & phi1)
			 | (OP==`ADC_izx & T==`Tthree & phi1)
			 | (OP==`ADC_izx & T==`Tfour & phi1)
			 | (OP==`ADC_izx & T==`Tfive & phi1)
			 | (OP==`ADC_zp & T==`Tzero & phi1)
			 | (OP==`ROR_zp & T==`Tzero & phi1)
			 | (OP==`ROR_zp & T==`Tthree & phi1)
			 | (OP==`ROR_zp & T==`Tfour & phi1)
			 | (OP==`PLA & T==`Tzero & phi1)
			 | (OP==`PLA & T==`Tthree & phi1)
			 | (OP==`JMP_zp & T==`Tzero & phi1)
			 | (OP==`JMP_zp & T==`Tfour & phi1)
			 | (OP==`ADC_abs & T==`Tzero & phi1)
			 | (OP==`ROR_abs & T==`Tzero & phi1)
			 | (OP==`ROR_abs & T==`Tfour & phi1)
			 | (OP==`ROR_abs & T==`Tfive & phi1)
			 | (OP==`ADC_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ADC_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`ADC_izy & T==`Tthree & phi1)
			 | (OP==`ADC_izy & T==`Tfour & phi1)
			 | (OP==`ADC_izy & T==`Tfive & phi1)
			 | (OP==`ADC_zpx & T==`Tzero & phi1)
			 | (OP==`ADC_zpx & T==`Tthree & phi1)
			 | (OP==`ROR_zpx & T==`Tzero & phi1)
			 | (OP==`ROR_zpx & T==`Tthree & phi1)
			 | (OP==`ROR_zpx & T==`Tfour & phi1)
			 | (OP==`ROR_zpx & T==`Tfive & phi1)
			 | (OP==`ADC_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ADC_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`ADC_aby & T==`Tfour & phi1)
			 | (OP==`ADC_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ADC_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`ADC_abx & T==`Tfour & phi1)
			 | (OP==`ROR_abx & T==`Tzero & phi1)
			 | (OP==`ROR_abx & T==`Tfour & phi1)
			 | (OP==`ROR_abx & T==`Tfive & phi1)
			 | (OP==`ROR_abx & T==`Tsix & phi1)
			 | (OP==`STA_izx & T==`Tzero & phi1)
			 | (OP==`STA_izx & T==`Tthree & phi1)
			 | (OP==`STA_izx & T==`Tfour & phi1)
			 | (OP==`STA_izx & T==`Tfive & phi1)
			 | (OP==`STY_zp & T==`Tzero & phi1)
			 | (OP==`STA_zp & T==`Tzero & phi1)
			 | (OP==`STX_zp & T==`Tzero & phi1)
			 | (OP==`STY_abs & T==`Tzero & phi1)
			 | (OP==`STA_abs & T==`Tzero & phi1)
			 | (OP==`STX_abs & T==`Tzero & phi1)
			 | (OP==`STA_izy & T==`Tzero & phi1)
			 | (OP==`STA_izy & T==`Tthree & phi1)
			 | (OP==`STA_izy & T==`Tfour & phi1)
			 | (OP==`STA_izy & T==`Tfive & phi1)
			 | (OP==`STY_zpx & T==`Tzero & phi1)
			 | (OP==`STY_zpx & T==`Tthree & phi1)
			 | (OP==`STA_zpx & T==`Tzero & phi1)
			 | (OP==`STA_zpx & T==`Tthree & phi1)
			 | (OP==`STX_zpy & T==`Tzero & phi1)
			 | (OP==`STX_zpy & T==`Tthree & phi1)
			 | (OP==`STA_aby & T==`Tzero & phi1)
			 | (OP==`STA_aby & T==`Tfour & phi1)
			 | (OP==`STA_abx & T==`Tzero & phi1)
			 | (OP==`STA_abx & T==`Tfour & phi1)
			 | (OP==`LDA_izx & T==`Tzero & phi1)
			 | (OP==`LDA_izx & T==`Tthree & phi1)
			 | (OP==`LDA_izx & T==`Tfour & phi1)
			 | (OP==`LDA_izx & T==`Tfive & phi1)
			 | (OP==`LDY_zp & T==`Tzero & phi1)
			 | (OP==`LDA_zp & T==`Tzero & phi1)
			 | (OP==`LDX_zp & T==`Tzero & phi1)
			 | (OP==`LDY_abs & T==`Tzero & phi1)
			 | (OP==`LDA_abs & T==`Tzero & phi1)
			 | (OP==`LDX_abs & T==`Tzero & phi1)
			 | (OP==`LDA_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDA_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`LDA_izy & T==`Tthree & phi1)
			 | (OP==`LDA_izy & T==`Tfour & phi1)
			 | (OP==`LDA_izy & T==`Tfive & phi1)
			 | (OP==`LDY_zpx & T==`Tzero & phi1)
			 | (OP==`LDY_zpx & T==`Tthree & phi1)
			 | (OP==`LDA_zpx & T==`Tzero & phi1)
			 | (OP==`LDA_zpx & T==`Tthree & phi1)
			 | (OP==`LDX_zpy & T==`Tzero & phi1)
			 | (OP==`LDX_zpy & T==`Tthree & phi1)
			 | (OP==`LDA_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDA_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`LDA_aby & T==`Tfour & phi1)
			 | (OP==`LDY_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDY_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`LDY_abx & T==`Tfour & phi1)
			 | (OP==`LDA_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDA_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`LDA_abx & T==`Tfour & phi1)
			 | (OP==`LDX_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDX_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`LDX_aby & T==`Tfour & phi1)
			 | (OP==`CMP_izx & T==`Tzero & phi1)
			 | (OP==`CMP_izx & T==`Tthree & phi1)
			 | (OP==`CMP_izx & T==`Tfour & phi1)
			 | (OP==`CMP_izx & T==`Tfive & phi1)
			 | (OP==`CPY_zp & T==`Tzero & phi1)
			 | (OP==`CMP_zp & T==`Tzero & phi1)
			 | (OP==`DEC_zp & T==`Tzero & phi1)
			 | (OP==`DEC_zp & T==`Tthree & phi1)
			 | (OP==`DEC_zp & T==`Tfour & phi1)
			 | (OP==`CPY_abs & T==`Tzero & phi1)
			 | (OP==`CMP_abs & T==`Tzero & phi1)
			 | (OP==`DEC_abs & T==`Tzero & phi1)
			 | (OP==`DEC_abs & T==`Tfour & phi1)
			 | (OP==`DEC_abs & T==`Tfive & phi1)
			 | (OP==`CMP_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`CMP_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`CMP_izy & T==`Tthree & phi1)
			 | (OP==`CMP_izy & T==`Tfour & phi1)
			 | (OP==`CMP_izy & T==`Tfive & phi1)
			 | (OP==`CMP_zpx & T==`Tzero & phi1)
			 | (OP==`CMP_zpx & T==`Tthree & phi1)
			 | (OP==`DEC_zpx & T==`Tzero & phi1)
			 | (OP==`DEC_zpx & T==`Tthree & phi1)
			 | (OP==`DEC_zpx & T==`Tfour & phi1)
			 | (OP==`DEC_zpx & T==`Tfive & phi1)
			 | (OP==`CMP_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`CMP_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`CMP_aby & T==`Tfour & phi1)
			 | (OP==`CMP_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`CMP_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`CMP_abx & T==`Tfour & phi1)
			 | (OP==`DEC_abx & T==`Tzero & phi1)
			 | (OP==`DEC_abx & T==`Tfour & phi1)
			 | (OP==`DEC_abx & T==`Tfive & phi1)
			 | (OP==`DEC_abx & T==`Tsix & phi1)
			 | (OP==`SBC_izx & T==`Tzero & phi1)
			 | (OP==`SBC_izx & T==`Tthree & phi1)
			 | (OP==`SBC_izx & T==`Tfour & phi1)
			 | (OP==`SBC_izx & T==`Tfive & phi1)
			 | (OP==`CPX_zp & T==`Tzero & phi1)
			 | (OP==`SBC_zp & T==`Tzero & phi1)
			 | (OP==`INC_zp & T==`Tzero & phi1)
			 | (OP==`INC_zp & T==`Tthree & phi1)
			 | (OP==`INC_zp & T==`Tfour & phi1)
			 | (OP==`CPX_abs & T==`Tzero & phi1)
			 | (OP==`SBC_abs & T==`Tzero & phi1)
			 | (OP==`INC_abs & T==`Tzero & phi1)
			 | (OP==`INC_abs & T==`Tfour & phi1)
			 | (OP==`INC_abs & T==`Tfive & phi1)
			 | (OP==`SBC_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`SBC_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`SBC_izy & T==`Tthree & phi1)
			 | (OP==`SBC_izy & T==`Tfour & phi1)
			 | (OP==`SBC_izy & T==`Tfive & phi1)
			 | (OP==`SBC_zpx & T==`Tzero & phi1)
			 | (OP==`SBC_zpx & T==`Tthree & phi1)
			 | (OP==`INC_zpx & T==`Tzero & phi1)
			 | (OP==`INC_zpx & T==`Tthree & phi1)
			 | (OP==`INC_zpx & T==`Tfour & phi1)
			 | (OP==`INC_zpx & T==`Tfive & phi1)
			 | (OP==`SBC_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`SBC_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`SBC_aby & T==`Tfour & phi1)
			 | (OP==`SBC_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`SBC_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`SBC_abx & T==`Tfour & phi1)
			 | (OP==`INC_abx & T==`Tzero & phi1)
			 | (OP==`INC_abx & T==`Tfour & phi1)
			 | (OP==`INC_abx & T==`Tfive & phi1)
			 | (OP==`INC_abx & T==`Tsix & phi1)
			;

assign control[`ADH_PCH] = (OP==`BRK & T==`Tone & phi1)
			 | (OP==`BRK & T==`Ttwo & phi1)
			 | (OP==`ORA_izx & T==`Tone & phi1)
			 | (OP==`ORA_izx & T==`Ttwo & phi1)
			 | (OP==`ORA_zp & T==`Tone & phi1)
			 | (OP==`ORA_zp & T==`Ttwo & phi1)
			 | (OP==`ASL_zp & T==`Tone & phi1)
			 | (OP==`ASL_zp & T==`Ttwo & phi1)
			 | (OP==`PHP & T==`Tone & phi1)
			 | (OP==`PHP & T==`Ttwo & phi1)
			 | (OP==`ORA_imm & T==`Tone & phi1)
			 | (OP==`ORA_imm & T==`Ttwo & phi1)
			 | (OP==`ASL & T==`Tone & phi1)
			 | (OP==`ASL & T==`Ttwo & phi1)
			 | (OP==`ORA_abs & T==`Tone & phi1)
			 | (OP==`ORA_abs & T==`Ttwo & phi1)
			 | (OP==`ORA_abs & T==`Tthree & phi1)
			 | (OP==`ASL_abs & T==`Tone & phi1)
			 | (OP==`ASL_abs & T==`Ttwo & phi1)
			 | (OP==`ASL_abs & T==`Tthree & phi1)
			 | (OP==`BPL_rel & T==`Tzero & phi1)
			 | (OP==`BPL_rel & T==`Ttwo & phi1)
			 | (OP==`BPL_rel & T==`Tthree & phi1)
			 | (OP==`BPL_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BPL_rel & T==`T1BranchCross & phi1)
			 | (OP==`BPL_rel & T==`T1NoBranch & phi1)
			 | (OP==`ORA_izy & T==`Tone & phi1)
			 | (OP==`ORA_izy & T==`Ttwo & phi1)
			 | (OP==`ORA_zpx & T==`Tone & phi1)
			 | (OP==`ORA_zpx & T==`Ttwo & phi1)
			 | (OP==`ASL_zpx & T==`Tone & phi1)
			 | (OP==`ASL_zpx & T==`Ttwo & phi1)
			 | (OP==`CLC & T==`Tone & phi1)
			 | (OP==`CLC & T==`Ttwo & phi1)
			 | (OP==`ORA_aby & T==`Tone & phi1)
			 | (OP==`ORA_aby & T==`Ttwo & phi1)
			 | (OP==`ORA_aby & T==`Tthree & phi1)
			 | (OP==`ORA_abx & T==`Tone & phi1)
			 | (OP==`ORA_abx & T==`Ttwo & phi1)
			 | (OP==`ORA_abx & T==`Tthree & phi1)
			 | (OP==`ASL_abx & T==`Tone & phi1)
			 | (OP==`ASL_abx & T==`Ttwo & phi1)
			 | (OP==`ASL_abx & T==`Tthree & phi1)
			 | (OP==`JSR_abs & T==`Tone & phi1)
			 | (OP==`JSR_abs & T==`Ttwo & phi1)
			 | (OP==`AND_izx & T==`Tone & phi1)
			 | (OP==`AND_izx & T==`Ttwo & phi1)
			 | (OP==`BIT_zp & T==`Tone & phi1)
			 | (OP==`BIT_zp & T==`Ttwo & phi1)
			 | (OP==`AND_zp & T==`Tone & phi1)
			 | (OP==`AND_zp & T==`Ttwo & phi1)
			 | (OP==`ROL_zp & T==`Tone & phi1)
			 | (OP==`ROL_zp & T==`Ttwo & phi1)
			 | (OP==`PLP & T==`Tone & phi1)
			 | (OP==`PLP & T==`Ttwo & phi1)
			 | (OP==`AND_imm & T==`Tone & phi1)
			 | (OP==`AND_imm & T==`Ttwo & phi1)
			 | (OP==`ROL & T==`Tone & phi1)
			 | (OP==`ROL & T==`Ttwo & phi1)
			 | (OP==`BIT_abs & T==`Tone & phi1)
			 | (OP==`BIT_abs & T==`Ttwo & phi1)
			 | (OP==`BIT_abs & T==`Tthree & phi1)
			 | (OP==`AND_abs & T==`Tone & phi1)
			 | (OP==`AND_abs & T==`Ttwo & phi1)
			 | (OP==`AND_abs & T==`Tthree & phi1)
			 | (OP==`ROL_abs & T==`Tone & phi1)
			 | (OP==`ROL_abs & T==`Ttwo & phi1)
			 | (OP==`ROL_abs & T==`Tthree & phi1)
			 | (OP==`BMI_rel & T==`Tzero & phi1)
			 | (OP==`BMI_rel & T==`Ttwo & phi1)
			 | (OP==`BMI_rel & T==`Tthree & phi1)
			 | (OP==`BMI_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BMI_rel & T==`T1BranchCross & phi1)
			 | (OP==`BMI_rel & T==`T1NoBranch & phi1)
			 | (OP==`AND_izy & T==`Tone & phi1)
			 | (OP==`AND_izy & T==`Ttwo & phi1)
			 | (OP==`AND_zpx & T==`Tone & phi1)
			 | (OP==`AND_zpx & T==`Ttwo & phi1)
			 | (OP==`ROL_zpx & T==`Tone & phi1)
			 | (OP==`ROL_zpx & T==`Ttwo & phi1)
			 | (OP==`SEC & T==`Tone & phi1)
			 | (OP==`SEC & T==`Ttwo & phi1)
			 | (OP==`AND_aby & T==`Tone & phi1)
			 | (OP==`AND_aby & T==`Ttwo & phi1)
			 | (OP==`AND_aby & T==`Tthree & phi1)
			 | (OP==`AND_abx & T==`Tone & phi1)
			 | (OP==`AND_abx & T==`Ttwo & phi1)
			 | (OP==`AND_abx & T==`Tthree & phi1)
			 | (OP==`ROL_abx & T==`Tone & phi1)
			 | (OP==`ROL_abx & T==`Ttwo & phi1)
			 | (OP==`ROL_abx & T==`Tthree & phi1)
			 | (OP==`RTI & T==`Tone & phi1)
			 | (OP==`RTI & T==`Ttwo & phi1)
			 | (OP==`EOR_izx & T==`Tone & phi1)
			 | (OP==`EOR_izx & T==`Ttwo & phi1)
			 | (OP==`EOR_zp & T==`Tone & phi1)
			 | (OP==`EOR_zp & T==`Ttwo & phi1)
			 | (OP==`LSR_zp & T==`Tone & phi1)
			 | (OP==`LSR_zp & T==`Ttwo & phi1)
			 | (OP==`PHA & T==`Tone & phi1)
			 | (OP==`PHA & T==`Ttwo & phi1)
			 | (OP==`EOR_imm & T==`Tone & phi1)
			 | (OP==`EOR_imm & T==`Ttwo & phi1)
			 | (OP==`LSR & T==`Tone & phi1)
			 | (OP==`LSR & T==`Ttwo & phi1)
			 | (OP==`JMP_abs & T==`Tzero & phi1)
			 | (OP==`JMP_abs & T==`Tone & phi1)
			 | (OP==`JMP_abs & T==`Ttwo & phi1)
			 | (OP==`EOR_abs & T==`Tone & phi1)
			 | (OP==`EOR_abs & T==`Ttwo & phi1)
			 | (OP==`EOR_abs & T==`Tthree & phi1)
			 | (OP==`LSR_abs & T==`Tone & phi1)
			 | (OP==`LSR_abs & T==`Ttwo & phi1)
			 | (OP==`LSR_abs & T==`Tthree & phi1)
			 | (OP==`BVC_rel & T==`Tzero & phi1)
			 | (OP==`BVC_rel & T==`Ttwo & phi1)
			 | (OP==`BVC_rel & T==`Tthree & phi1)
			 | (OP==`BVC_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BVC_rel & T==`T1BranchCross & phi1)
			 | (OP==`BVC_rel & T==`T1NoBranch & phi1)
			 | (OP==`EOR_izy & T==`Tone & phi1)
			 | (OP==`EOR_izy & T==`Ttwo & phi1)
			 | (OP==`EOR_zpx & T==`Tone & phi1)
			 | (OP==`EOR_zpx & T==`Ttwo & phi1)
			 | (OP==`LSR_zpx & T==`Tone & phi1)
			 | (OP==`LSR_zpx & T==`Ttwo & phi1)
			 | (OP==`CLI & T==`Tone & phi1)
			 | (OP==`CLI & T==`Ttwo & phi1)
			 | (OP==`EOR_aby & T==`Tone & phi1)
			 | (OP==`EOR_aby & T==`Ttwo & phi1)
			 | (OP==`EOR_aby & T==`Tthree & phi1)
			 | (OP==`EOR_abx & T==`Tone & phi1)
			 | (OP==`EOR_abx & T==`Ttwo & phi1)
			 | (OP==`EOR_abx & T==`Tthree & phi1)
			 | (OP==`LSR_abx & T==`Tone & phi1)
			 | (OP==`LSR_abx & T==`Ttwo & phi1)
			 | (OP==`LSR_abx & T==`Tthree & phi1)
			 | (OP==`RTS & T==`Tzero & phi1)
			 | (OP==`RTS & T==`Tone & phi1)
			 | (OP==`RTS & T==`Ttwo & phi1)
			 | (OP==`ADC_izx & T==`Tone & phi1)
			 | (OP==`ADC_izx & T==`Ttwo & phi1)
			 | (OP==`ADC_zp & T==`Tone & phi1)
			 | (OP==`ADC_zp & T==`Ttwo & phi1)
			 | (OP==`ROR_zp & T==`Tone & phi1)
			 | (OP==`ROR_zp & T==`Ttwo & phi1)
			 | (OP==`PLA & T==`Tone & phi1)
			 | (OP==`PLA & T==`Ttwo & phi1)
			 | (OP==`ADC_imm & T==`Tone & phi1)
			 | (OP==`ADC_imm & T==`Ttwo & phi1)
			 | (OP==`ROR & T==`Tone & phi1)
			 | (OP==`ROR & T==`Ttwo & phi1)
			 | (OP==`JMP_zp & T==`Tone & phi1)
			 | (OP==`JMP_zp & T==`Ttwo & phi1)
			 | (OP==`JMP_zp & T==`Tthree & phi1)
			 | (OP==`ADC_abs & T==`Tone & phi1)
			 | (OP==`ADC_abs & T==`Ttwo & phi1)
			 | (OP==`ADC_abs & T==`Tthree & phi1)
			 | (OP==`ROR_abs & T==`Tone & phi1)
			 | (OP==`ROR_abs & T==`Ttwo & phi1)
			 | (OP==`ROR_abs & T==`Tthree & phi1)
			 | (OP==`BVS_rel & T==`Tzero & phi1)
			 | (OP==`BVS_rel & T==`Ttwo & phi1)
			 | (OP==`BVS_rel & T==`Tthree & phi1)
			 | (OP==`BVS_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BVS_rel & T==`T1BranchCross & phi1)
			 | (OP==`BVS_rel & T==`T1NoBranch & phi1)
			 | (OP==`ADC_izy & T==`Tone & phi1)
			 | (OP==`ADC_izy & T==`Ttwo & phi1)
			 | (OP==`ADC_zpx & T==`Tone & phi1)
			 | (OP==`ADC_zpx & T==`Ttwo & phi1)
			 | (OP==`ROR_zpx & T==`Tone & phi1)
			 | (OP==`ROR_zpx & T==`Ttwo & phi1)
			 | (OP==`SEI & T==`Tone & phi1)
			 | (OP==`SEI & T==`Ttwo & phi1)
			 | (OP==`ADC_aby & T==`Tone & phi1)
			 | (OP==`ADC_aby & T==`Ttwo & phi1)
			 | (OP==`ADC_aby & T==`Tthree & phi1)
			 | (OP==`ADC_abx & T==`Tone & phi1)
			 | (OP==`ADC_abx & T==`Ttwo & phi1)
			 | (OP==`ADC_abx & T==`Tthree & phi1)
			 | (OP==`ROR_abx & T==`Tone & phi1)
			 | (OP==`ROR_abx & T==`Ttwo & phi1)
			 | (OP==`ROR_abx & T==`Tthree & phi1)
			 | (OP==`STA_izx & T==`Tone & phi1)
			 | (OP==`STA_izx & T==`Ttwo & phi1)
			 | (OP==`STY_zp & T==`Tone & phi1)
			 | (OP==`STY_zp & T==`Ttwo & phi1)
			 | (OP==`STA_zp & T==`Tone & phi1)
			 | (OP==`STA_zp & T==`Ttwo & phi1)
			 | (OP==`STX_zp & T==`Tone & phi1)
			 | (OP==`STX_zp & T==`Ttwo & phi1)
			 | (OP==`DEY & T==`Tone & phi1)
			 | (OP==`DEY & T==`Ttwo & phi1)
			 | (OP==`TXA & T==`Tone & phi1)
			 | (OP==`TXA & T==`Ttwo & phi1)
			 | (OP==`STY_abs & T==`Tone & phi1)
			 | (OP==`STY_abs & T==`Ttwo & phi1)
			 | (OP==`STY_abs & T==`Tthree & phi1)
			 | (OP==`STA_abs & T==`Tone & phi1)
			 | (OP==`STA_abs & T==`Ttwo & phi1)
			 | (OP==`STA_abs & T==`Tthree & phi1)
			 | (OP==`STX_abs & T==`Tone & phi1)
			 | (OP==`STX_abs & T==`Ttwo & phi1)
			 | (OP==`STX_abs & T==`Tthree & phi1)
			 | (OP==`BCC_rel & T==`Tzero & phi1)
			 | (OP==`BCC_rel & T==`Ttwo & phi1)
			 | (OP==`BCC_rel & T==`Tthree & phi1)
			 | (OP==`BCC_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BCC_rel & T==`T1BranchCross & phi1)
			 | (OP==`BCC_rel & T==`T1NoBranch & phi1)
			 | (OP==`STA_izy & T==`Tone & phi1)
			 | (OP==`STA_izy & T==`Ttwo & phi1)
			 | (OP==`STY_zpx & T==`Tone & phi1)
			 | (OP==`STY_zpx & T==`Ttwo & phi1)
			 | (OP==`STA_zpx & T==`Tone & phi1)
			 | (OP==`STA_zpx & T==`Ttwo & phi1)
			 | (OP==`STX_zpy & T==`Tone & phi1)
			 | (OP==`STX_zpy & T==`Ttwo & phi1)
			 | (OP==`TYA & T==`Tone & phi1)
			 | (OP==`TYA & T==`Ttwo & phi1)
			 | (OP==`STA_aby & T==`Tone & phi1)
			 | (OP==`STA_aby & T==`Ttwo & phi1)
			 | (OP==`STA_aby & T==`Tthree & phi1)
			 | (OP==`TXS & T==`Tone & phi1)
			 | (OP==`TXS & T==`Ttwo & phi1)
			 | (OP==`STA_abx & T==`Tone & phi1)
			 | (OP==`STA_abx & T==`Ttwo & phi1)
			 | (OP==`STA_abx & T==`Tthree & phi1)
			 | (OP==`LDY_imm & T==`Tone & phi1)
			 | (OP==`LDY_imm & T==`Ttwo & phi1)
			 | (OP==`LDA_izx & T==`Tone & phi1)
			 | (OP==`LDA_izx & T==`Ttwo & phi1)
			 | (OP==`LDX_imm & T==`Tone & phi1)
			 | (OP==`LDX_imm & T==`Ttwo & phi1)
			 | (OP==`LDY_zp & T==`Tone & phi1)
			 | (OP==`LDY_zp & T==`Ttwo & phi1)
			 | (OP==`LDA_zp & T==`Tone & phi1)
			 | (OP==`LDA_zp & T==`Ttwo & phi1)
			 | (OP==`LDX_zp & T==`Tone & phi1)
			 | (OP==`LDX_zp & T==`Ttwo & phi1)
			 | (OP==`TAY & T==`Tone & phi1)
			 | (OP==`TAY & T==`Ttwo & phi1)
			 | (OP==`LDA_imm & T==`Tone & phi1)
			 | (OP==`LDA_imm & T==`Ttwo & phi1)
			 | (OP==`TAX & T==`Tone & phi1)
			 | (OP==`TAX & T==`Ttwo & phi1)
			 | (OP==`LDY_abs & T==`Tone & phi1)
			 | (OP==`LDY_abs & T==`Ttwo & phi1)
			 | (OP==`LDY_abs & T==`Tthree & phi1)
			 | (OP==`LDA_abs & T==`Tone & phi1)
			 | (OP==`LDA_abs & T==`Ttwo & phi1)
			 | (OP==`LDA_abs & T==`Tthree & phi1)
			 | (OP==`LDX_abs & T==`Tone & phi1)
			 | (OP==`LDX_abs & T==`Ttwo & phi1)
			 | (OP==`LDX_abs & T==`Tthree & phi1)
			 | (OP==`BCS_rel & T==`Tzero & phi1)
			 | (OP==`BCS_rel & T==`Ttwo & phi1)
			 | (OP==`BCS_rel & T==`Tthree & phi1)
			 | (OP==`BCS_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BCS_rel & T==`T1BranchCross & phi1)
			 | (OP==`BCS_rel & T==`T1NoBranch & phi1)
			 | (OP==`LDA_izy & T==`Tone & phi1)
			 | (OP==`LDA_izy & T==`Ttwo & phi1)
			 | (OP==`LDY_zpx & T==`Tone & phi1)
			 | (OP==`LDY_zpx & T==`Ttwo & phi1)
			 | (OP==`LDA_zpx & T==`Tone & phi1)
			 | (OP==`LDA_zpx & T==`Ttwo & phi1)
			 | (OP==`LDX_zpy & T==`Tone & phi1)
			 | (OP==`LDX_zpy & T==`Ttwo & phi1)
			 | (OP==`CLV & T==`Tone & phi1)
			 | (OP==`CLV & T==`Ttwo & phi1)
			 | (OP==`LDA_aby & T==`Tone & phi1)
			 | (OP==`LDA_aby & T==`Ttwo & phi1)
			 | (OP==`LDA_aby & T==`Tthree & phi1)
			 | (OP==`TSX & T==`Tone & phi1)
			 | (OP==`TSX & T==`Ttwo & phi1)
			 | (OP==`LDY_abx & T==`Tone & phi1)
			 | (OP==`LDY_abx & T==`Ttwo & phi1)
			 | (OP==`LDY_abx & T==`Tthree & phi1)
			 | (OP==`LDA_abx & T==`Tone & phi1)
			 | (OP==`LDA_abx & T==`Ttwo & phi1)
			 | (OP==`LDA_abx & T==`Tthree & phi1)
			 | (OP==`LDX_aby & T==`Tone & phi1)
			 | (OP==`LDX_aby & T==`Ttwo & phi1)
			 | (OP==`LDX_aby & T==`Tthree & phi1)
			 | (OP==`CPY_imm & T==`Tone & phi1)
			 | (OP==`CPY_imm & T==`Ttwo & phi1)
			 | (OP==`CMP_izx & T==`Tone & phi1)
			 | (OP==`CMP_izx & T==`Ttwo & phi1)
			 | (OP==`CPY_zp & T==`Tone & phi1)
			 | (OP==`CPY_zp & T==`Ttwo & phi1)
			 | (OP==`CMP_zp & T==`Tone & phi1)
			 | (OP==`CMP_zp & T==`Ttwo & phi1)
			 | (OP==`DEC_zp & T==`Tone & phi1)
			 | (OP==`DEC_zp & T==`Ttwo & phi1)
			 | (OP==`INY & T==`Tone & phi1)
			 | (OP==`INY & T==`Ttwo & phi1)
			 | (OP==`CMP_imm & T==`Tone & phi1)
			 | (OP==`CMP_imm & T==`Ttwo & phi1)
			 | (OP==`DEX & T==`Tone & phi1)
			 | (OP==`DEX & T==`Ttwo & phi1)
			 | (OP==`CPY_abs & T==`Tone & phi1)
			 | (OP==`CPY_abs & T==`Ttwo & phi1)
			 | (OP==`CPY_abs & T==`Tthree & phi1)
			 | (OP==`CMP_abs & T==`Tone & phi1)
			 | (OP==`CMP_abs & T==`Ttwo & phi1)
			 | (OP==`CMP_abs & T==`Tthree & phi1)
			 | (OP==`DEC_abs & T==`Tone & phi1)
			 | (OP==`DEC_abs & T==`Ttwo & phi1)
			 | (OP==`DEC_abs & T==`Tthree & phi1)
			 | (OP==`BNE_rel & T==`Tzero & phi1)
			 | (OP==`BNE_rel & T==`Ttwo & phi1)
			 | (OP==`BNE_rel & T==`Tthree & phi1)
			 | (OP==`BNE_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BNE_rel & T==`T1BranchCross & phi1)
			 | (OP==`BNE_rel & T==`T1NoBranch & phi1)
			 | (OP==`CMP_izy & T==`Tone & phi1)
			 | (OP==`CMP_izy & T==`Ttwo & phi1)
			 | (OP==`CMP_zpx & T==`Tone & phi1)
			 | (OP==`CMP_zpx & T==`Ttwo & phi1)
			 | (OP==`DEC_zpx & T==`Tone & phi1)
			 | (OP==`DEC_zpx & T==`Ttwo & phi1)
			 | (OP==`CLD & T==`Tone & phi1)
			 | (OP==`CLD & T==`Ttwo & phi1)
			 | (OP==`CMP_aby & T==`Tone & phi1)
			 | (OP==`CMP_aby & T==`Ttwo & phi1)
			 | (OP==`CMP_aby & T==`Tthree & phi1)
			 | (OP==`CMP_abx & T==`Tone & phi1)
			 | (OP==`CMP_abx & T==`Ttwo & phi1)
			 | (OP==`CMP_abx & T==`Tthree & phi1)
			 | (OP==`DEC_abx & T==`Tone & phi1)
			 | (OP==`DEC_abx & T==`Ttwo & phi1)
			 | (OP==`DEC_abx & T==`Tthree & phi1)
			 | (OP==`CPX_imm & T==`Tone & phi1)
			 | (OP==`CPX_imm & T==`Ttwo & phi1)
			 | (OP==`SBC_izx & T==`Tone & phi1)
			 | (OP==`SBC_izx & T==`Ttwo & phi1)
			 | (OP==`CPX_zp & T==`Tone & phi1)
			 | (OP==`CPX_zp & T==`Ttwo & phi1)
			 | (OP==`SBC_zp & T==`Tone & phi1)
			 | (OP==`SBC_zp & T==`Ttwo & phi1)
			 | (OP==`INC_zp & T==`Tone & phi1)
			 | (OP==`INC_zp & T==`Ttwo & phi1)
			 | (OP==`INX & T==`Tone & phi1)
			 | (OP==`INX & T==`Ttwo & phi1)
			 | (OP==`SBC_imm & T==`Tone & phi1)
			 | (OP==`SBC_imm & T==`Ttwo & phi1)
			 | (OP==`NOP & T==`Tone & phi1)
			 | (OP==`NOP & T==`Ttwo & phi1)
			 | (OP==`CPX_abs & T==`Tone & phi1)
			 | (OP==`CPX_abs & T==`Ttwo & phi1)
			 | (OP==`CPX_abs & T==`Tthree & phi1)
			 | (OP==`SBC_abs & T==`Tone & phi1)
			 | (OP==`SBC_abs & T==`Ttwo & phi1)
			 | (OP==`SBC_abs & T==`Tthree & phi1)
			 | (OP==`INC_abs & T==`Tone & phi1)
			 | (OP==`INC_abs & T==`Ttwo & phi1)
			 | (OP==`INC_abs & T==`Tthree & phi1)
			 | (OP==`BEQ_rel & T==`Tzero & phi1)
			 | (OP==`BEQ_rel & T==`Ttwo & phi1)
			 | (OP==`BEQ_rel & T==`Tthree & phi1)
			 | (OP==`BEQ_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BEQ_rel & T==`T1BranchCross & phi1)
			 | (OP==`BEQ_rel & T==`T1NoBranch & phi1)
			 | (OP==`SBC_izy & T==`Tone & phi1)
			 | (OP==`SBC_izy & T==`Ttwo & phi1)
			 | (OP==`SBC_zpx & T==`Tone & phi1)
			 | (OP==`SBC_zpx & T==`Ttwo & phi1)
			 | (OP==`INC_zpx & T==`Tone & phi1)
			 | (OP==`INC_zpx & T==`Ttwo & phi1)
			 | (OP==`SED & T==`Tone & phi1)
			 | (OP==`SED & T==`Ttwo & phi1)
			 | (OP==`SBC_aby & T==`Tone & phi1)
			 | (OP==`SBC_aby & T==`Ttwo & phi1)
			 | (OP==`SBC_aby & T==`Tthree & phi1)
			 | (OP==`SBC_abx & T==`Tone & phi1)
			 | (OP==`SBC_abx & T==`Ttwo & phi1)
			 | (OP==`SBC_abx & T==`Tthree & phi1)
			 | (OP==`INC_abx & T==`Tone & phi1)
			 | (OP==`INC_abx & T==`Ttwo & phi1)
			 | (OP==`INC_abx & T==`Tthree & phi1)
			;

assign control[`PCH_DB] = (OP==`BRK & T==`Ttwo & phi2)
			 | (OP==`BRK & T==`Tthree & phi1)
			 | (OP==`JSR_abs & T==`Tthree & phi2)
			 | (OP==`JSR_abs & T==`Tfour & phi1)
			;

assign control[`PCH_ADH] = (OP==`BRK & T==`Tone & phi2)
			 | (OP==`BRK & T==`Ttwo & phi1)
			 | (OP==`ORA_izx & T==`Tzero & phi2)
			 | (OP==`ORA_izx & T==`Tone & phi1)
			 | (OP==`ORA_izx & T==`Tone & phi2)
			 | (OP==`ORA_izx & T==`Ttwo & phi1)
			 | (OP==`ORA_zp & T==`Tzero & phi2)
			 | (OP==`ORA_zp & T==`Tone & phi1)
			 | (OP==`ORA_zp & T==`Tone & phi2)
			 | (OP==`ORA_zp & T==`Ttwo & phi1)
			 | (OP==`ASL_zp & T==`Tzero & phi2)
			 | (OP==`ASL_zp & T==`Tone & phi1)
			 | (OP==`ASL_zp & T==`Tone & phi2)
			 | (OP==`ASL_zp & T==`Ttwo & phi1)
			 | (OP==`PHP & T==`Tzero & phi2)
			 | (OP==`PHP & T==`Tone & phi1)
			 | (OP==`PHP & T==`Tone & phi2)
			 | (OP==`PHP & T==`Ttwo & phi1)
			 | (OP==`ORA_imm & T==`Tone & phi1)
			 | (OP==`ORA_imm & T==`Tone & phi2)
			 | (OP==`ORA_imm & T==`Ttwo & phi1)
			 | (OP==`ORA_imm & T==`Ttwo & phi2)
			 | (OP==`ASL & T==`Tone & phi1)
			 | (OP==`ASL & T==`Tone & phi2)
			 | (OP==`ASL & T==`Ttwo & phi1)
			 | (OP==`ASL & T==`Ttwo & phi2)
			 | (OP==`ORA_abs & T==`Tzero & phi2)
			 | (OP==`ORA_abs & T==`Tone & phi1)
			 | (OP==`ORA_abs & T==`Tone & phi2)
			 | (OP==`ORA_abs & T==`Ttwo & phi1)
			 | (OP==`ORA_abs & T==`Ttwo & phi2)
			 | (OP==`ORA_abs & T==`Tthree & phi1)
			 | (OP==`ASL_abs & T==`Tzero & phi2)
			 | (OP==`ASL_abs & T==`Tone & phi1)
			 | (OP==`ASL_abs & T==`Tone & phi2)
			 | (OP==`ASL_abs & T==`Ttwo & phi1)
			 | (OP==`ASL_abs & T==`Ttwo & phi2)
			 | (OP==`ASL_abs & T==`Tthree & phi1)
			 | (OP==`BPL_rel & T==`Tzero & phi1)
			 | (OP==`BPL_rel & T==`Ttwo & phi1)
			 | (OP==`BPL_rel & T==`Ttwo & phi2)
			 | (OP==`BPL_rel & T==`Tthree & phi1)
			 | (OP==`BPL_rel & T==`Tthree & phi2)
			 | (OP==`BPL_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BPL_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BPL_rel & T==`T1BranchCross & phi2)
			 | (OP==`BPL_rel & T==`T1NoBranch & phi1)
			 | (OP==`BPL_rel & T==`T1NoBranch & phi2)
			 | (OP==`ORA_izy & T==`TzeroCrossPg & phi2)
			 | (OP==`ORA_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`ORA_izy & T==`Tone & phi1)
			 | (OP==`ORA_izy & T==`Tone & phi2)
			 | (OP==`ORA_izy & T==`Ttwo & phi1)
			 | (OP==`ORA_zpx & T==`Tzero & phi2)
			 | (OP==`ORA_zpx & T==`Tone & phi1)
			 | (OP==`ORA_zpx & T==`Tone & phi2)
			 | (OP==`ORA_zpx & T==`Ttwo & phi1)
			 | (OP==`ASL_zpx & T==`Tzero & phi2)
			 | (OP==`ASL_zpx & T==`Tone & phi1)
			 | (OP==`ASL_zpx & T==`Tone & phi2)
			 | (OP==`ASL_zpx & T==`Ttwo & phi1)
			 | (OP==`CLC & T==`Tone & phi1)
			 | (OP==`CLC & T==`Tone & phi2)
			 | (OP==`CLC & T==`Ttwo & phi1)
			 | (OP==`CLC & T==`Ttwo & phi2)
			 | (OP==`ORA_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`ORA_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`ORA_aby & T==`Tone & phi1)
			 | (OP==`ORA_aby & T==`Tone & phi2)
			 | (OP==`ORA_aby & T==`Ttwo & phi1)
			 | (OP==`ORA_aby & T==`Ttwo & phi2)
			 | (OP==`ORA_aby & T==`Tthree & phi1)
			 | (OP==`ORA_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`ORA_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`ORA_abx & T==`Tone & phi1)
			 | (OP==`ORA_abx & T==`Tone & phi2)
			 | (OP==`ORA_abx & T==`Ttwo & phi1)
			 | (OP==`ORA_abx & T==`Ttwo & phi2)
			 | (OP==`ORA_abx & T==`Tthree & phi1)
			 | (OP==`ASL_abx & T==`Tzero & phi2)
			 | (OP==`ASL_abx & T==`Tone & phi1)
			 | (OP==`ASL_abx & T==`Tone & phi2)
			 | (OP==`ASL_abx & T==`Ttwo & phi1)
			 | (OP==`ASL_abx & T==`Ttwo & phi2)
			 | (OP==`ASL_abx & T==`Tthree & phi1)
			 | (OP==`JSR_abs & T==`Tzero & phi1)
			 | (OP==`JSR_abs & T==`Tone & phi2)
			 | (OP==`JSR_abs & T==`Ttwo & phi1)
			 | (OP==`JSR_abs & T==`Tfive & phi2)
			 | (OP==`AND_izx & T==`Tzero & phi2)
			 | (OP==`AND_izx & T==`Tone & phi1)
			 | (OP==`AND_izx & T==`Tone & phi2)
			 | (OP==`AND_izx & T==`Ttwo & phi1)
			 | (OP==`BIT_zp & T==`Tzero & phi2)
			 | (OP==`BIT_zp & T==`Tone & phi1)
			 | (OP==`BIT_zp & T==`Tone & phi2)
			 | (OP==`BIT_zp & T==`Ttwo & phi1)
			 | (OP==`AND_zp & T==`Tzero & phi2)
			 | (OP==`AND_zp & T==`Tone & phi1)
			 | (OP==`AND_zp & T==`Tone & phi2)
			 | (OP==`AND_zp & T==`Ttwo & phi1)
			 | (OP==`ROL_zp & T==`Tzero & phi2)
			 | (OP==`ROL_zp & T==`Tone & phi1)
			 | (OP==`ROL_zp & T==`Tone & phi2)
			 | (OP==`ROL_zp & T==`Ttwo & phi1)
			 | (OP==`PLP & T==`Tzero & phi2)
			 | (OP==`PLP & T==`Tone & phi1)
			 | (OP==`PLP & T==`Tone & phi2)
			 | (OP==`PLP & T==`Ttwo & phi1)
			 | (OP==`AND_imm & T==`Tone & phi1)
			 | (OP==`AND_imm & T==`Tone & phi2)
			 | (OP==`AND_imm & T==`Ttwo & phi1)
			 | (OP==`AND_imm & T==`Ttwo & phi2)
			 | (OP==`ROL & T==`Tone & phi1)
			 | (OP==`ROL & T==`Tone & phi2)
			 | (OP==`ROL & T==`Ttwo & phi1)
			 | (OP==`ROL & T==`Ttwo & phi2)
			 | (OP==`BIT_abs & T==`Tzero & phi2)
			 | (OP==`BIT_abs & T==`Tone & phi1)
			 | (OP==`BIT_abs & T==`Tone & phi2)
			 | (OP==`BIT_abs & T==`Ttwo & phi1)
			 | (OP==`BIT_abs & T==`Ttwo & phi2)
			 | (OP==`BIT_abs & T==`Tthree & phi1)
			 | (OP==`AND_abs & T==`Tzero & phi2)
			 | (OP==`AND_abs & T==`Tone & phi1)
			 | (OP==`AND_abs & T==`Tone & phi2)
			 | (OP==`AND_abs & T==`Ttwo & phi1)
			 | (OP==`AND_abs & T==`Ttwo & phi2)
			 | (OP==`AND_abs & T==`Tthree & phi1)
			 | (OP==`ROL_abs & T==`Tzero & phi2)
			 | (OP==`ROL_abs & T==`Tone & phi1)
			 | (OP==`ROL_abs & T==`Tone & phi2)
			 | (OP==`ROL_abs & T==`Ttwo & phi1)
			 | (OP==`ROL_abs & T==`Ttwo & phi2)
			 | (OP==`ROL_abs & T==`Tthree & phi1)
			 | (OP==`BMI_rel & T==`Tzero & phi1)
			 | (OP==`BMI_rel & T==`Ttwo & phi1)
			 | (OP==`BMI_rel & T==`Ttwo & phi2)
			 | (OP==`BMI_rel & T==`Tthree & phi1)
			 | (OP==`BMI_rel & T==`Tthree & phi2)
			 | (OP==`BMI_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BMI_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BMI_rel & T==`T1BranchCross & phi2)
			 | (OP==`BMI_rel & T==`T1NoBranch & phi1)
			 | (OP==`BMI_rel & T==`T1NoBranch & phi2)
			 | (OP==`AND_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`AND_izy & T==`TzeroCrossPg & phi2)
			 | (OP==`AND_izy & T==`Tone & phi1)
			 | (OP==`AND_izy & T==`Tone & phi2)
			 | (OP==`AND_izy & T==`Ttwo & phi1)
			 | (OP==`AND_zpx & T==`Tzero & phi2)
			 | (OP==`AND_zpx & T==`Tone & phi1)
			 | (OP==`AND_zpx & T==`Tone & phi2)
			 | (OP==`AND_zpx & T==`Ttwo & phi1)
			 | (OP==`ROL_zpx & T==`Tzero & phi2)
			 | (OP==`ROL_zpx & T==`Tone & phi1)
			 | (OP==`ROL_zpx & T==`Tone & phi2)
			 | (OP==`ROL_zpx & T==`Ttwo & phi1)
			 | (OP==`SEC & T==`Tone & phi1)
			 | (OP==`SEC & T==`Tone & phi2)
			 | (OP==`SEC & T==`Ttwo & phi1)
			 | (OP==`SEC & T==`Ttwo & phi2)
			 | (OP==`AND_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`AND_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`AND_aby & T==`Tone & phi1)
			 | (OP==`AND_aby & T==`Tone & phi2)
			 | (OP==`AND_aby & T==`Ttwo & phi1)
			 | (OP==`AND_aby & T==`Ttwo & phi2)
			 | (OP==`AND_aby & T==`Tthree & phi1)
			 | (OP==`AND_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`AND_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`AND_abx & T==`Tone & phi1)
			 | (OP==`AND_abx & T==`Tone & phi2)
			 | (OP==`AND_abx & T==`Ttwo & phi1)
			 | (OP==`AND_abx & T==`Ttwo & phi2)
			 | (OP==`AND_abx & T==`Tthree & phi1)
			 | (OP==`ROL_abx & T==`Tzero & phi2)
			 | (OP==`ROL_abx & T==`Tone & phi1)
			 | (OP==`ROL_abx & T==`Tone & phi2)
			 | (OP==`ROL_abx & T==`Ttwo & phi1)
			 | (OP==`ROL_abx & T==`Ttwo & phi2)
			 | (OP==`ROL_abx & T==`Tthree & phi1)
			 | (OP==`RTI & T==`Tone & phi2)
			 | (OP==`RTI & T==`Ttwo & phi1)
			 | (OP==`EOR_izx & T==`Tzero & phi2)
			 | (OP==`EOR_izx & T==`Tone & phi1)
			 | (OP==`EOR_izx & T==`Tone & phi2)
			 | (OP==`EOR_izx & T==`Ttwo & phi1)
			 | (OP==`EOR_zp & T==`Tzero & phi2)
			 | (OP==`EOR_zp & T==`Tone & phi1)
			 | (OP==`EOR_zp & T==`Tone & phi2)
			 | (OP==`EOR_zp & T==`Ttwo & phi1)
			 | (OP==`LSR_zp & T==`Tzero & phi2)
			 | (OP==`LSR_zp & T==`Tone & phi1)
			 | (OP==`LSR_zp & T==`Tone & phi2)
			 | (OP==`LSR_zp & T==`Ttwo & phi1)
			 | (OP==`PHA & T==`Tzero & phi2)
			 | (OP==`PHA & T==`Tone & phi1)
			 | (OP==`PHA & T==`Tone & phi2)
			 | (OP==`PHA & T==`Ttwo & phi1)
			 | (OP==`EOR_imm & T==`Tone & phi1)
			 | (OP==`EOR_imm & T==`Tone & phi2)
			 | (OP==`EOR_imm & T==`Ttwo & phi1)
			 | (OP==`EOR_imm & T==`Ttwo & phi2)
			 | (OP==`LSR & T==`Tone & phi1)
			 | (OP==`LSR & T==`Tone & phi2)
			 | (OP==`LSR & T==`Ttwo & phi1)
			 | (OP==`LSR & T==`Ttwo & phi2)
			 | (OP==`JMP_abs & T==`Tzero & phi1)
			 | (OP==`JMP_abs & T==`Tone & phi2)
			 | (OP==`JMP_abs & T==`Ttwo & phi1)
			 | (OP==`JMP_abs & T==`Ttwo & phi2)
			 | (OP==`EOR_abs & T==`Tzero & phi2)
			 | (OP==`EOR_abs & T==`Tone & phi1)
			 | (OP==`EOR_abs & T==`Tone & phi2)
			 | (OP==`EOR_abs & T==`Ttwo & phi1)
			 | (OP==`EOR_abs & T==`Ttwo & phi2)
			 | (OP==`EOR_abs & T==`Tthree & phi1)
			 | (OP==`LSR_abs & T==`Tzero & phi2)
			 | (OP==`LSR_abs & T==`Tone & phi1)
			 | (OP==`LSR_abs & T==`Tone & phi2)
			 | (OP==`LSR_abs & T==`Ttwo & phi1)
			 | (OP==`LSR_abs & T==`Ttwo & phi2)
			 | (OP==`LSR_abs & T==`Tthree & phi1)
			 | (OP==`BVC_rel & T==`Tzero & phi1)
			 | (OP==`BVC_rel & T==`Ttwo & phi1)
			 | (OP==`BVC_rel & T==`Ttwo & phi2)
			 | (OP==`BVC_rel & T==`Tthree & phi1)
			 | (OP==`BVC_rel & T==`Tthree & phi2)
			 | (OP==`BVC_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BVC_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BVC_rel & T==`T1BranchCross & phi2)
			 | (OP==`BVC_rel & T==`T1NoBranch & phi1)
			 | (OP==`BVC_rel & T==`T1NoBranch & phi2)
			 | (OP==`EOR_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`EOR_izy & T==`TzeroCrossPg & phi2)
			 | (OP==`EOR_izy & T==`Tone & phi1)
			 | (OP==`EOR_izy & T==`Tone & phi2)
			 | (OP==`EOR_izy & T==`Ttwo & phi1)
			 | (OP==`EOR_zpx & T==`Tzero & phi2)
			 | (OP==`EOR_zpx & T==`Tone & phi1)
			 | (OP==`EOR_zpx & T==`Tone & phi2)
			 | (OP==`EOR_zpx & T==`Ttwo & phi1)
			 | (OP==`LSR_zpx & T==`Tzero & phi2)
			 | (OP==`LSR_zpx & T==`Tone & phi1)
			 | (OP==`LSR_zpx & T==`Tone & phi2)
			 | (OP==`LSR_zpx & T==`Ttwo & phi1)
			 | (OP==`CLI & T==`Tone & phi1)
			 | (OP==`CLI & T==`Tone & phi2)
			 | (OP==`CLI & T==`Ttwo & phi1)
			 | (OP==`CLI & T==`Ttwo & phi2)
			 | (OP==`EOR_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`EOR_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`EOR_aby & T==`Tone & phi1)
			 | (OP==`EOR_aby & T==`Tone & phi2)
			 | (OP==`EOR_aby & T==`Ttwo & phi1)
			 | (OP==`EOR_aby & T==`Ttwo & phi2)
			 | (OP==`EOR_aby & T==`Tthree & phi1)
			 | (OP==`EOR_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`EOR_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`EOR_abx & T==`Tone & phi1)
			 | (OP==`EOR_abx & T==`Tone & phi2)
			 | (OP==`EOR_abx & T==`Ttwo & phi1)
			 | (OP==`EOR_abx & T==`Ttwo & phi2)
			 | (OP==`EOR_abx & T==`Tthree & phi1)
			 | (OP==`LSR_abx & T==`Tzero & phi2)
			 | (OP==`LSR_abx & T==`Tone & phi1)
			 | (OP==`LSR_abx & T==`Tone & phi2)
			 | (OP==`LSR_abx & T==`Ttwo & phi1)
			 | (OP==`LSR_abx & T==`Ttwo & phi2)
			 | (OP==`LSR_abx & T==`Tthree & phi1)
			 | (OP==`RTS & T==`Tzero & phi2)
			 | (OP==`RTS & T==`Tone & phi1)
			 | (OP==`RTS & T==`Tone & phi2)
			 | (OP==`RTS & T==`Ttwo & phi1)
			 | (OP==`ADC_izx & T==`Tzero & phi2)
			 | (OP==`ADC_izx & T==`Tone & phi1)
			 | (OP==`ADC_izx & T==`Tone & phi2)
			 | (OP==`ADC_izx & T==`Ttwo & phi1)
			 | (OP==`ADC_zp & T==`Tzero & phi2)
			 | (OP==`ADC_zp & T==`Tone & phi1)
			 | (OP==`ADC_zp & T==`Tone & phi2)
			 | (OP==`ADC_zp & T==`Ttwo & phi1)
			 | (OP==`ROR_zp & T==`Tzero & phi2)
			 | (OP==`ROR_zp & T==`Tone & phi1)
			 | (OP==`ROR_zp & T==`Tone & phi2)
			 | (OP==`ROR_zp & T==`Ttwo & phi1)
			 | (OP==`PLA & T==`Tzero & phi2)
			 | (OP==`PLA & T==`Tone & phi1)
			 | (OP==`PLA & T==`Tone & phi2)
			 | (OP==`PLA & T==`Ttwo & phi1)
			 | (OP==`ADC_imm & T==`Tone & phi1)
			 | (OP==`ADC_imm & T==`Tone & phi2)
			 | (OP==`ADC_imm & T==`Ttwo & phi1)
			 | (OP==`ADC_imm & T==`Ttwo & phi2)
			 | (OP==`ROR & T==`Tone & phi1)
			 | (OP==`ROR & T==`Tone & phi2)
			 | (OP==`ROR & T==`Ttwo & phi1)
			 | (OP==`ROR & T==`Ttwo & phi2)
			 | (OP==`JMP_zp & T==`Tone & phi2)
			 | (OP==`JMP_zp & T==`Ttwo & phi1)
			 | (OP==`JMP_zp & T==`Ttwo & phi2)
			 | (OP==`JMP_zp & T==`Tthree & phi1)
			 | (OP==`ADC_abs & T==`Tzero & phi2)
			 | (OP==`ADC_abs & T==`Tone & phi1)
			 | (OP==`ADC_abs & T==`Tone & phi2)
			 | (OP==`ADC_abs & T==`Ttwo & phi1)
			 | (OP==`ADC_abs & T==`Ttwo & phi2)
			 | (OP==`ADC_abs & T==`Tthree & phi1)
			 | (OP==`ROR_abs & T==`Tzero & phi2)
			 | (OP==`ROR_abs & T==`Tone & phi1)
			 | (OP==`ROR_abs & T==`Tone & phi2)
			 | (OP==`ROR_abs & T==`Ttwo & phi1)
			 | (OP==`ROR_abs & T==`Ttwo & phi2)
			 | (OP==`ROR_abs & T==`Tthree & phi1)
			 | (OP==`BVS_rel & T==`Tzero & phi1)
			 | (OP==`BVS_rel & T==`Ttwo & phi1)
			 | (OP==`BVS_rel & T==`Ttwo & phi2)
			 | (OP==`BVS_rel & T==`Tthree & phi1)
			 | (OP==`BVS_rel & T==`Tthree & phi2)
			 | (OP==`BVS_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BVS_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BVS_rel & T==`T1BranchCross & phi2)
			 | (OP==`BVS_rel & T==`T1NoBranch & phi1)
			 | (OP==`BVS_rel & T==`T1NoBranch & phi2)
			 | (OP==`ADC_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`ADC_izy & T==`TzeroCrossPg & phi2)
			 | (OP==`ADC_izy & T==`Tone & phi1)
			 | (OP==`ADC_izy & T==`Tone & phi2)
			 | (OP==`ADC_izy & T==`Ttwo & phi1)
			 | (OP==`ADC_zpx & T==`Tzero & phi2)
			 | (OP==`ADC_zpx & T==`Tone & phi1)
			 | (OP==`ADC_zpx & T==`Tone & phi2)
			 | (OP==`ADC_zpx & T==`Ttwo & phi1)
			 | (OP==`ROR_zpx & T==`Tzero & phi2)
			 | (OP==`ROR_zpx & T==`Tone & phi1)
			 | (OP==`ROR_zpx & T==`Tone & phi2)
			 | (OP==`ROR_zpx & T==`Ttwo & phi1)
			 | (OP==`SEI & T==`Tone & phi1)
			 | (OP==`SEI & T==`Tone & phi2)
			 | (OP==`SEI & T==`Ttwo & phi1)
			 | (OP==`SEI & T==`Ttwo & phi2)
			 | (OP==`ADC_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`ADC_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`ADC_aby & T==`Tone & phi1)
			 | (OP==`ADC_aby & T==`Tone & phi2)
			 | (OP==`ADC_aby & T==`Ttwo & phi1)
			 | (OP==`ADC_aby & T==`Ttwo & phi2)
			 | (OP==`ADC_aby & T==`Tthree & phi1)
			 | (OP==`ADC_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`ADC_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`ADC_abx & T==`Tone & phi1)
			 | (OP==`ADC_abx & T==`Tone & phi2)
			 | (OP==`ADC_abx & T==`Ttwo & phi1)
			 | (OP==`ADC_abx & T==`Ttwo & phi2)
			 | (OP==`ADC_abx & T==`Tthree & phi1)
			 | (OP==`ROR_abx & T==`Tzero & phi2)
			 | (OP==`ROR_abx & T==`Tone & phi1)
			 | (OP==`ROR_abx & T==`Tone & phi2)
			 | (OP==`ROR_abx & T==`Ttwo & phi1)
			 | (OP==`ROR_abx & T==`Ttwo & phi2)
			 | (OP==`ROR_abx & T==`Tthree & phi1)
			 | (OP==`STA_izx & T==`Tzero & phi2)
			 | (OP==`STA_izx & T==`Tone & phi1)
			 | (OP==`STA_izx & T==`Tone & phi2)
			 | (OP==`STA_izx & T==`Ttwo & phi1)
			 | (OP==`STY_zp & T==`Tzero & phi2)
			 | (OP==`STY_zp & T==`Tone & phi1)
			 | (OP==`STY_zp & T==`Tone & phi2)
			 | (OP==`STY_zp & T==`Ttwo & phi1)
			 | (OP==`STA_zp & T==`Tzero & phi2)
			 | (OP==`STA_zp & T==`Tone & phi1)
			 | (OP==`STA_zp & T==`Tone & phi2)
			 | (OP==`STA_zp & T==`Ttwo & phi1)
			 | (OP==`STX_zp & T==`Tzero & phi2)
			 | (OP==`STX_zp & T==`Tone & phi1)
			 | (OP==`STX_zp & T==`Tone & phi2)
			 | (OP==`STX_zp & T==`Ttwo & phi1)
			 | (OP==`DEY & T==`Tone & phi1)
			 | (OP==`DEY & T==`Tone & phi2)
			 | (OP==`DEY & T==`Ttwo & phi1)
			 | (OP==`DEY & T==`Ttwo & phi2)
			 | (OP==`TXA & T==`Tone & phi1)
			 | (OP==`TXA & T==`Tone & phi2)
			 | (OP==`TXA & T==`Ttwo & phi1)
			 | (OP==`TXA & T==`Ttwo & phi2)
			 | (OP==`STY_abs & T==`Tzero & phi2)
			 | (OP==`STY_abs & T==`Tone & phi1)
			 | (OP==`STY_abs & T==`Tone & phi2)
			 | (OP==`STY_abs & T==`Ttwo & phi1)
			 | (OP==`STY_abs & T==`Ttwo & phi2)
			 | (OP==`STY_abs & T==`Tthree & phi1)
			 | (OP==`STA_abs & T==`Tzero & phi2)
			 | (OP==`STA_abs & T==`Tone & phi1)
			 | (OP==`STA_abs & T==`Tone & phi2)
			 | (OP==`STA_abs & T==`Ttwo & phi1)
			 | (OP==`STA_abs & T==`Ttwo & phi2)
			 | (OP==`STA_abs & T==`Tthree & phi1)
			 | (OP==`STX_abs & T==`Tzero & phi2)
			 | (OP==`STX_abs & T==`Tone & phi1)
			 | (OP==`STX_abs & T==`Tone & phi2)
			 | (OP==`STX_abs & T==`Ttwo & phi1)
			 | (OP==`STX_abs & T==`Ttwo & phi2)
			 | (OP==`STX_abs & T==`Tthree & phi1)
			 | (OP==`BCC_rel & T==`Tzero & phi1)
			 | (OP==`BCC_rel & T==`Ttwo & phi1)
			 | (OP==`BCC_rel & T==`Ttwo & phi2)
			 | (OP==`BCC_rel & T==`Tthree & phi1)
			 | (OP==`BCC_rel & T==`Tthree & phi2)
			 | (OP==`BCC_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BCC_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BCC_rel & T==`T1BranchCross & phi2)
			 | (OP==`BCC_rel & T==`T1NoBranch & phi1)
			 | (OP==`BCC_rel & T==`T1NoBranch & phi2)
			 | (OP==`STA_izy & T==`Tzero & phi2)
			 | (OP==`STA_izy & T==`Tone & phi1)
			 | (OP==`STA_izy & T==`Tone & phi2)
			 | (OP==`STA_izy & T==`Ttwo & phi1)
			 | (OP==`STY_zpx & T==`Tzero & phi2)
			 | (OP==`STY_zpx & T==`Tone & phi1)
			 | (OP==`STY_zpx & T==`Tone & phi2)
			 | (OP==`STY_zpx & T==`Ttwo & phi1)
			 | (OP==`STA_zpx & T==`Tzero & phi2)
			 | (OP==`STA_zpx & T==`Tone & phi1)
			 | (OP==`STA_zpx & T==`Tone & phi2)
			 | (OP==`STA_zpx & T==`Ttwo & phi1)
			 | (OP==`STX_zpy & T==`Tzero & phi2)
			 | (OP==`STX_zpy & T==`Tone & phi1)
			 | (OP==`STX_zpy & T==`Tone & phi2)
			 | (OP==`STX_zpy & T==`Ttwo & phi1)
			 | (OP==`TYA & T==`Tone & phi1)
			 | (OP==`TYA & T==`Tone & phi2)
			 | (OP==`TYA & T==`Ttwo & phi1)
			 | (OP==`TYA & T==`Ttwo & phi2)
			 | (OP==`STA_aby & T==`Tzero & phi2)
			 | (OP==`STA_aby & T==`Tone & phi1)
			 | (OP==`STA_aby & T==`Tone & phi2)
			 | (OP==`STA_aby & T==`Ttwo & phi1)
			 | (OP==`STA_aby & T==`Ttwo & phi2)
			 | (OP==`STA_aby & T==`Tthree & phi1)
			 | (OP==`TXS & T==`Tone & phi1)
			 | (OP==`TXS & T==`Tone & phi2)
			 | (OP==`TXS & T==`Ttwo & phi1)
			 | (OP==`TXS & T==`Ttwo & phi2)
			 | (OP==`STA_abx & T==`Tzero & phi2)
			 | (OP==`STA_abx & T==`Tone & phi1)
			 | (OP==`STA_abx & T==`Tone & phi2)
			 | (OP==`STA_abx & T==`Ttwo & phi1)
			 | (OP==`STA_abx & T==`Ttwo & phi2)
			 | (OP==`STA_abx & T==`Tthree & phi1)
			 | (OP==`LDY_imm & T==`Tone & phi1)
			 | (OP==`LDY_imm & T==`Tone & phi2)
			 | (OP==`LDY_imm & T==`Ttwo & phi1)
			 | (OP==`LDY_imm & T==`Ttwo & phi2)
			 | (OP==`LDA_izx & T==`Tzero & phi2)
			 | (OP==`LDA_izx & T==`Tone & phi1)
			 | (OP==`LDA_izx & T==`Tone & phi2)
			 | (OP==`LDA_izx & T==`Ttwo & phi1)
			 | (OP==`LDX_imm & T==`Tone & phi1)
			 | (OP==`LDX_imm & T==`Tone & phi2)
			 | (OP==`LDX_imm & T==`Ttwo & phi1)
			 | (OP==`LDX_imm & T==`Ttwo & phi2)
			 | (OP==`LDY_zp & T==`Tzero & phi2)
			 | (OP==`LDY_zp & T==`Tone & phi1)
			 | (OP==`LDY_zp & T==`Tone & phi2)
			 | (OP==`LDY_zp & T==`Ttwo & phi1)
			 | (OP==`LDA_zp & T==`Tzero & phi2)
			 | (OP==`LDA_zp & T==`Tone & phi1)
			 | (OP==`LDA_zp & T==`Tone & phi2)
			 | (OP==`LDA_zp & T==`Ttwo & phi1)
			 | (OP==`LDX_zp & T==`Tzero & phi2)
			 | (OP==`LDX_zp & T==`Tone & phi1)
			 | (OP==`LDX_zp & T==`Tone & phi2)
			 | (OP==`LDX_zp & T==`Ttwo & phi1)
			 | (OP==`TAY & T==`Tone & phi1)
			 | (OP==`TAY & T==`Tone & phi2)
			 | (OP==`TAY & T==`Ttwo & phi1)
			 | (OP==`TAY & T==`Ttwo & phi2)
			 | (OP==`LDA_imm & T==`Tone & phi1)
			 | (OP==`LDA_imm & T==`Tone & phi2)
			 | (OP==`LDA_imm & T==`Ttwo & phi1)
			 | (OP==`LDA_imm & T==`Ttwo & phi2)
			 | (OP==`TAX & T==`Tone & phi1)
			 | (OP==`TAX & T==`Tone & phi2)
			 | (OP==`TAX & T==`Ttwo & phi1)
			 | (OP==`TAX & T==`Ttwo & phi2)
			 | (OP==`LDY_abs & T==`Tzero & phi2)
			 | (OP==`LDY_abs & T==`Tone & phi1)
			 | (OP==`LDY_abs & T==`Tone & phi2)
			 | (OP==`LDY_abs & T==`Ttwo & phi1)
			 | (OP==`LDY_abs & T==`Ttwo & phi2)
			 | (OP==`LDY_abs & T==`Tthree & phi1)
			 | (OP==`LDA_abs & T==`Tzero & phi2)
			 | (OP==`LDA_abs & T==`Tone & phi1)
			 | (OP==`LDA_abs & T==`Tone & phi2)
			 | (OP==`LDA_abs & T==`Ttwo & phi1)
			 | (OP==`LDA_abs & T==`Ttwo & phi2)
			 | (OP==`LDA_abs & T==`Tthree & phi1)
			 | (OP==`LDX_abs & T==`Tzero & phi2)
			 | (OP==`LDX_abs & T==`Tone & phi1)
			 | (OP==`LDX_abs & T==`Tone & phi2)
			 | (OP==`LDX_abs & T==`Ttwo & phi1)
			 | (OP==`LDX_abs & T==`Ttwo & phi2)
			 | (OP==`LDX_abs & T==`Tthree & phi1)
			 | (OP==`BCS_rel & T==`Tzero & phi1)
			 | (OP==`BCS_rel & T==`Ttwo & phi1)
			 | (OP==`BCS_rel & T==`Ttwo & phi2)
			 | (OP==`BCS_rel & T==`Tthree & phi1)
			 | (OP==`BCS_rel & T==`Tthree & phi2)
			 | (OP==`BCS_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BCS_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BCS_rel & T==`T1BranchCross & phi2)
			 | (OP==`BCS_rel & T==`T1NoBranch & phi1)
			 | (OP==`BCS_rel & T==`T1NoBranch & phi2)
			 | (OP==`LDA_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`LDA_izy & T==`TzeroCrossPg & phi2)
			 | (OP==`LDA_izy & T==`Tone & phi1)
			 | (OP==`LDA_izy & T==`Tone & phi2)
			 | (OP==`LDA_izy & T==`Ttwo & phi1)
			 | (OP==`LDY_zpx & T==`Tzero & phi2)
			 | (OP==`LDY_zpx & T==`Tone & phi1)
			 | (OP==`LDY_zpx & T==`Tone & phi2)
			 | (OP==`LDY_zpx & T==`Ttwo & phi1)
			 | (OP==`LDA_zpx & T==`Tzero & phi2)
			 | (OP==`LDA_zpx & T==`Tone & phi1)
			 | (OP==`LDA_zpx & T==`Tone & phi2)
			 | (OP==`LDA_zpx & T==`Ttwo & phi1)
			 | (OP==`LDX_zpy & T==`Tzero & phi2)
			 | (OP==`LDX_zpy & T==`Tone & phi1)
			 | (OP==`LDX_zpy & T==`Tone & phi2)
			 | (OP==`LDX_zpy & T==`Ttwo & phi1)
			 | (OP==`CLV & T==`Tone & phi1)
			 | (OP==`CLV & T==`Tone & phi2)
			 | (OP==`CLV & T==`Ttwo & phi1)
			 | (OP==`CLV & T==`Ttwo & phi2)
			 | (OP==`LDA_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`LDA_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`LDA_aby & T==`Tone & phi1)
			 | (OP==`LDA_aby & T==`Tone & phi2)
			 | (OP==`LDA_aby & T==`Ttwo & phi1)
			 | (OP==`LDA_aby & T==`Ttwo & phi2)
			 | (OP==`LDA_aby & T==`Tthree & phi1)
			 | (OP==`TSX & T==`Tone & phi1)
			 | (OP==`TSX & T==`Tone & phi2)
			 | (OP==`TSX & T==`Ttwo & phi1)
			 | (OP==`TSX & T==`Ttwo & phi2)
			 | (OP==`LDY_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`LDY_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`LDY_abx & T==`Tone & phi1)
			 | (OP==`LDY_abx & T==`Tone & phi2)
			 | (OP==`LDY_abx & T==`Ttwo & phi1)
			 | (OP==`LDY_abx & T==`Ttwo & phi2)
			 | (OP==`LDY_abx & T==`Tthree & phi1)
			 | (OP==`LDA_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`LDA_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`LDA_abx & T==`Tone & phi1)
			 | (OP==`LDA_abx & T==`Tone & phi2)
			 | (OP==`LDA_abx & T==`Ttwo & phi1)
			 | (OP==`LDA_abx & T==`Ttwo & phi2)
			 | (OP==`LDA_abx & T==`Tthree & phi1)
			 | (OP==`LDX_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`LDX_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`LDX_aby & T==`Tone & phi1)
			 | (OP==`LDX_aby & T==`Tone & phi2)
			 | (OP==`LDX_aby & T==`Ttwo & phi1)
			 | (OP==`LDX_aby & T==`Ttwo & phi2)
			 | (OP==`LDX_aby & T==`Tthree & phi1)
			 | (OP==`CPY_imm & T==`Tone & phi1)
			 | (OP==`CPY_imm & T==`Tone & phi2)
			 | (OP==`CPY_imm & T==`Ttwo & phi1)
			 | (OP==`CPY_imm & T==`Ttwo & phi2)
			 | (OP==`CMP_izx & T==`Tzero & phi2)
			 | (OP==`CMP_izx & T==`Tone & phi1)
			 | (OP==`CMP_izx & T==`Tone & phi2)
			 | (OP==`CMP_izx & T==`Ttwo & phi1)
			 | (OP==`CPY_zp & T==`Tzero & phi2)
			 | (OP==`CPY_zp & T==`Tone & phi1)
			 | (OP==`CPY_zp & T==`Tone & phi2)
			 | (OP==`CPY_zp & T==`Ttwo & phi1)
			 | (OP==`CMP_zp & T==`Tzero & phi2)
			 | (OP==`CMP_zp & T==`Tone & phi1)
			 | (OP==`CMP_zp & T==`Tone & phi2)
			 | (OP==`CMP_zp & T==`Ttwo & phi1)
			 | (OP==`DEC_zp & T==`Tzero & phi2)
			 | (OP==`DEC_zp & T==`Tone & phi1)
			 | (OP==`DEC_zp & T==`Tone & phi2)
			 | (OP==`DEC_zp & T==`Ttwo & phi1)
			 | (OP==`INY & T==`Tone & phi1)
			 | (OP==`INY & T==`Tone & phi2)
			 | (OP==`INY & T==`Ttwo & phi1)
			 | (OP==`INY & T==`Ttwo & phi2)
			 | (OP==`CMP_imm & T==`Tone & phi1)
			 | (OP==`CMP_imm & T==`Tone & phi2)
			 | (OP==`CMP_imm & T==`Ttwo & phi1)
			 | (OP==`CMP_imm & T==`Ttwo & phi2)
			 | (OP==`DEX & T==`Tone & phi1)
			 | (OP==`DEX & T==`Tone & phi2)
			 | (OP==`DEX & T==`Ttwo & phi1)
			 | (OP==`DEX & T==`Ttwo & phi2)
			 | (OP==`CPY_abs & T==`Tzero & phi2)
			 | (OP==`CPY_abs & T==`Tone & phi1)
			 | (OP==`CPY_abs & T==`Tone & phi2)
			 | (OP==`CPY_abs & T==`Ttwo & phi1)
			 | (OP==`CPY_abs & T==`Ttwo & phi2)
			 | (OP==`CPY_abs & T==`Tthree & phi1)
			 | (OP==`CMP_abs & T==`Tzero & phi2)
			 | (OP==`CMP_abs & T==`Tone & phi1)
			 | (OP==`CMP_abs & T==`Tone & phi2)
			 | (OP==`CMP_abs & T==`Ttwo & phi1)
			 | (OP==`CMP_abs & T==`Ttwo & phi2)
			 | (OP==`CMP_abs & T==`Tthree & phi1)
			 | (OP==`DEC_abs & T==`Tzero & phi2)
			 | (OP==`DEC_abs & T==`Tone & phi1)
			 | (OP==`DEC_abs & T==`Tone & phi2)
			 | (OP==`DEC_abs & T==`Ttwo & phi1)
			 | (OP==`DEC_abs & T==`Ttwo & phi2)
			 | (OP==`DEC_abs & T==`Tthree & phi1)
			 | (OP==`BNE_rel & T==`Tzero & phi1)
			 | (OP==`BNE_rel & T==`Ttwo & phi1)
			 | (OP==`BNE_rel & T==`Ttwo & phi2)
			 | (OP==`BNE_rel & T==`Tthree & phi1)
			 | (OP==`BNE_rel & T==`Tthree & phi2)
			 | (OP==`BNE_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BNE_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BNE_rel & T==`T1BranchCross & phi2)
			 | (OP==`BNE_rel & T==`T1NoBranch & phi1)
			 | (OP==`BNE_rel & T==`T1NoBranch & phi2)
			 | (OP==`CMP_izy & T==`TzeroCrossPg & phi2)
			 | (OP==`CMP_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`CMP_izy & T==`Tone & phi1)
			 | (OP==`CMP_izy & T==`Tone & phi2)
			 | (OP==`CMP_izy & T==`Ttwo & phi1)
			 | (OP==`CMP_zpx & T==`Tzero & phi2)
			 | (OP==`CMP_zpx & T==`Tone & phi1)
			 | (OP==`CMP_zpx & T==`Tone & phi2)
			 | (OP==`CMP_zpx & T==`Ttwo & phi1)
			 | (OP==`DEC_zpx & T==`Tzero & phi2)
			 | (OP==`DEC_zpx & T==`Tone & phi1)
			 | (OP==`DEC_zpx & T==`Tone & phi2)
			 | (OP==`DEC_zpx & T==`Ttwo & phi1)
			 | (OP==`CLD & T==`Tone & phi1)
			 | (OP==`CLD & T==`Tone & phi2)
			 | (OP==`CLD & T==`Ttwo & phi1)
			 | (OP==`CLD & T==`Ttwo & phi2)
			 | (OP==`CMP_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`CMP_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`CMP_aby & T==`Tone & phi1)
			 | (OP==`CMP_aby & T==`Tone & phi2)
			 | (OP==`CMP_aby & T==`Ttwo & phi1)
			 | (OP==`CMP_aby & T==`Ttwo & phi2)
			 | (OP==`CMP_aby & T==`Tthree & phi1)
			 | (OP==`CMP_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`CMP_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`CMP_abx & T==`Tone & phi1)
			 | (OP==`CMP_abx & T==`Tone & phi2)
			 | (OP==`CMP_abx & T==`Ttwo & phi1)
			 | (OP==`CMP_abx & T==`Ttwo & phi2)
			 | (OP==`CMP_abx & T==`Tthree & phi1)
			 | (OP==`DEC_abx & T==`Tzero & phi2)
			 | (OP==`DEC_abx & T==`Tone & phi1)
			 | (OP==`DEC_abx & T==`Tone & phi2)
			 | (OP==`DEC_abx & T==`Ttwo & phi1)
			 | (OP==`DEC_abx & T==`Ttwo & phi2)
			 | (OP==`DEC_abx & T==`Tthree & phi1)
			 | (OP==`CPX_imm & T==`Tone & phi1)
			 | (OP==`CPX_imm & T==`Tone & phi2)
			 | (OP==`CPX_imm & T==`Ttwo & phi1)
			 | (OP==`CPX_imm & T==`Ttwo & phi2)
			 | (OP==`SBC_izx & T==`Tzero & phi2)
			 | (OP==`SBC_izx & T==`Tone & phi1)
			 | (OP==`SBC_izx & T==`Tone & phi2)
			 | (OP==`SBC_izx & T==`Ttwo & phi1)
			 | (OP==`CPX_zp & T==`Tzero & phi2)
			 | (OP==`CPX_zp & T==`Tone & phi1)
			 | (OP==`CPX_zp & T==`Tone & phi2)
			 | (OP==`CPX_zp & T==`Ttwo & phi1)
			 | (OP==`SBC_zp & T==`Tzero & phi2)
			 | (OP==`SBC_zp & T==`Tone & phi1)
			 | (OP==`SBC_zp & T==`Tone & phi2)
			 | (OP==`SBC_zp & T==`Ttwo & phi1)
			 | (OP==`INC_zp & T==`Tzero & phi2)
			 | (OP==`INC_zp & T==`Tone & phi1)
			 | (OP==`INC_zp & T==`Tone & phi2)
			 | (OP==`INC_zp & T==`Ttwo & phi1)
			 | (OP==`INX & T==`Tone & phi1)
			 | (OP==`INX & T==`Tone & phi2)
			 | (OP==`INX & T==`Ttwo & phi1)
			 | (OP==`INX & T==`Ttwo & phi2)
			 | (OP==`SBC_imm & T==`Tone & phi1)
			 | (OP==`SBC_imm & T==`Tone & phi2)
			 | (OP==`SBC_imm & T==`Ttwo & phi1)
			 | (OP==`SBC_imm & T==`Ttwo & phi2)
			 | (OP==`NOP & T==`Tone & phi1)
			 | (OP==`NOP & T==`Tone & phi2)
			 | (OP==`NOP & T==`Ttwo & phi1)
			 | (OP==`NOP & T==`Ttwo & phi2)
			 | (OP==`CPX_abs & T==`Tzero & phi2)
			 | (OP==`CPX_abs & T==`Tone & phi1)
			 | (OP==`CPX_abs & T==`Tone & phi2)
			 | (OP==`CPX_abs & T==`Ttwo & phi1)
			 | (OP==`CPX_abs & T==`Ttwo & phi2)
			 | (OP==`CPX_abs & T==`Tthree & phi1)
			 | (OP==`SBC_abs & T==`Tzero & phi2)
			 | (OP==`SBC_abs & T==`Tone & phi1)
			 | (OP==`SBC_abs & T==`Tone & phi2)
			 | (OP==`SBC_abs & T==`Ttwo & phi1)
			 | (OP==`SBC_abs & T==`Ttwo & phi2)
			 | (OP==`SBC_abs & T==`Tthree & phi1)
			 | (OP==`INC_abs & T==`Tzero & phi2)
			 | (OP==`INC_abs & T==`Tone & phi1)
			 | (OP==`INC_abs & T==`Tone & phi2)
			 | (OP==`INC_abs & T==`Ttwo & phi1)
			 | (OP==`INC_abs & T==`Ttwo & phi2)
			 | (OP==`INC_abs & T==`Tthree & phi1)
			 | (OP==`BEQ_rel & T==`Tzero & phi1)
			 | (OP==`BEQ_rel & T==`Ttwo & phi1)
			 | (OP==`BEQ_rel & T==`Ttwo & phi2)
			 | (OP==`BEQ_rel & T==`Tthree & phi1)
			 | (OP==`BEQ_rel & T==`Tthree & phi2)
			 | (OP==`BEQ_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BEQ_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BEQ_rel & T==`T1BranchCross & phi2)
			 | (OP==`BEQ_rel & T==`T1NoBranch & phi1)
			 | (OP==`BEQ_rel & T==`T1NoBranch & phi2)
			 | (OP==`SBC_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`SBC_izy & T==`TzeroCrossPg & phi2)
			 | (OP==`SBC_izy & T==`Tone & phi1)
			 | (OP==`SBC_izy & T==`Tone & phi2)
			 | (OP==`SBC_izy & T==`Ttwo & phi1)
			 | (OP==`SBC_zpx & T==`Tzero & phi2)
			 | (OP==`SBC_zpx & T==`Tone & phi1)
			 | (OP==`SBC_zpx & T==`Tone & phi2)
			 | (OP==`SBC_zpx & T==`Ttwo & phi1)
			 | (OP==`INC_zpx & T==`Tzero & phi2)
			 | (OP==`INC_zpx & T==`Tone & phi1)
			 | (OP==`INC_zpx & T==`Tone & phi2)
			 | (OP==`INC_zpx & T==`Ttwo & phi1)
			 | (OP==`SED & T==`Tone & phi1)
			 | (OP==`SED & T==`Tone & phi2)
			 | (OP==`SED & T==`Ttwo & phi1)
			 | (OP==`SED & T==`Ttwo & phi2)
			 | (OP==`SBC_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`SBC_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`SBC_aby & T==`Tone & phi1)
			 | (OP==`SBC_aby & T==`Tone & phi2)
			 | (OP==`SBC_aby & T==`Ttwo & phi1)
			 | (OP==`SBC_aby & T==`Ttwo & phi2)
			 | (OP==`SBC_aby & T==`Tthree & phi1)
			 | (OP==`SBC_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`SBC_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`SBC_abx & T==`Tone & phi1)
			 | (OP==`SBC_abx & T==`Tone & phi2)
			 | (OP==`SBC_abx & T==`Ttwo & phi1)
			 | (OP==`SBC_abx & T==`Ttwo & phi2)
			 | (OP==`SBC_abx & T==`Tthree & phi1)
			 | (OP==`INC_abx & T==`Tzero & phi2)
			 | (OP==`INC_abx & T==`Tone & phi1)
			 | (OP==`INC_abx & T==`Tone & phi2)
			 | (OP==`INC_abx & T==`Ttwo & phi1)
			 | (OP==`INC_abx & T==`Ttwo & phi2)
			 | (OP==`INC_abx & T==`Tthree & phi1)
			;

assign control[`SB_ADH] = (OP==`BPL_rel & T==`Tzero & phi1)
			 | (OP==`BPL_rel & T==`Tzero & phi2)
			 | (OP==`BPL_rel & T==`Tthree & phi2)
			 | (OP==`BPL_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BPL_rel & T==`T1BranchCross & phi1)
			 | (OP==`ORA_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`ORA_izy & T==`Tfive & phi2)
			 | (OP==`ORA_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`ORA_aby & T==`Tfour & phi2)
			 | (OP==`ORA_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`ORA_abx & T==`Tfour & phi2)
			 | (OP==`ASL_abx & T==`Tfour & phi2)
			 | (OP==`ASL_abx & T==`Tfive & phi1)
			 | (OP==`BMI_rel & T==`Tzero & phi1)
			 | (OP==`BMI_rel & T==`Tzero & phi2)
			 | (OP==`BMI_rel & T==`Tthree & phi2)
			 | (OP==`BMI_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BMI_rel & T==`T1BranchCross & phi1)
			 | (OP==`AND_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`AND_izy & T==`Tfive & phi2)
			 | (OP==`AND_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`AND_aby & T==`Tfour & phi2)
			 | (OP==`AND_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`AND_abx & T==`Tfour & phi2)
			 | (OP==`ROL_abx & T==`Tfour & phi2)
			 | (OP==`ROL_abx & T==`Tfive & phi1)
			 | (OP==`BVC_rel & T==`Tzero & phi1)
			 | (OP==`BVC_rel & T==`Tzero & phi2)
			 | (OP==`BVC_rel & T==`Tthree & phi2)
			 | (OP==`BVC_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BVC_rel & T==`T1BranchCross & phi1)
			 | (OP==`EOR_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`EOR_izy & T==`Tfive & phi2)
			 | (OP==`EOR_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`EOR_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`EOR_aby & T==`Tfour & phi2)
			 | (OP==`EOR_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`EOR_abx & T==`Tfour & phi2)
			 | (OP==`LSR_abx & T==`Tfour & phi2)
			 | (OP==`LSR_abx & T==`Tfive & phi1)
			 | (OP==`BVS_rel & T==`Tzero & phi1)
			 | (OP==`BVS_rel & T==`Tzero & phi2)
			 | (OP==`BVS_rel & T==`Tthree & phi2)
			 | (OP==`BVS_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BVS_rel & T==`T1BranchCross & phi1)
			 | (OP==`ADC_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`ADC_izy & T==`Tfive & phi2)
			 | (OP==`ADC_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`ADC_aby & T==`Tfour & phi2)
			 | (OP==`ADC_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`ADC_abx & T==`Tfour & phi2)
			 | (OP==`ROR_abx & T==`Tfour & phi2)
			 | (OP==`ROR_abx & T==`Tfive & phi1)
			 | (OP==`BCC_rel & T==`Tzero & phi1)
			 | (OP==`BCC_rel & T==`Tzero & phi2)
			 | (OP==`BCC_rel & T==`Tthree & phi2)
			 | (OP==`BCC_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BCC_rel & T==`T1BranchCross & phi1)
			 | (OP==`STA_izy & T==`Tzero & phi1)
			 | (OP==`STA_izy & T==`Tfive & phi2)
			 | (OP==`STA_aby & T==`Tzero & phi1)
			 | (OP==`STA_aby & T==`Tfour & phi2)
			 | (OP==`STA_abx & T==`Tzero & phi1)
			 | (OP==`STA_abx & T==`Tfour & phi2)
			 | (OP==`BCS_rel & T==`Tzero & phi1)
			 | (OP==`BCS_rel & T==`Tzero & phi2)
			 | (OP==`BCS_rel & T==`Tthree & phi2)
			 | (OP==`BCS_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BCS_rel & T==`T1BranchCross & phi1)
			 | (OP==`LDA_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`LDA_izy & T==`Tfive & phi2)
			 | (OP==`LDA_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`LDA_aby & T==`Tfour & phi2)
			 | (OP==`LDY_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`LDY_abx & T==`Tfour & phi2)
			 | (OP==`LDA_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`LDA_abx & T==`Tfour & phi2)
			 | (OP==`LDX_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`LDX_aby & T==`Tfour & phi2)
			 | (OP==`BNE_rel & T==`Tzero & phi1)
			 | (OP==`BNE_rel & T==`Tzero & phi2)
			 | (OP==`BNE_rel & T==`Tthree & phi2)
			 | (OP==`BNE_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BNE_rel & T==`T1BranchCross & phi1)
			 | (OP==`CMP_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`CMP_izy & T==`Tfive & phi2)
			 | (OP==`CMP_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`CMP_aby & T==`Tfour & phi2)
			 | (OP==`CMP_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`CMP_abx & T==`Tfour & phi2)
			 | (OP==`DEC_abx & T==`Tfour & phi2)
			 | (OP==`DEC_abx & T==`Tfive & phi1)
			 | (OP==`BEQ_rel & T==`Tzero & phi1)
			 | (OP==`BEQ_rel & T==`Tzero & phi2)
			 | (OP==`BEQ_rel & T==`Tthree & phi2)
			 | (OP==`BEQ_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BEQ_rel & T==`T1BranchCross & phi1)
			 | (OP==`SBC_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`SBC_izy & T==`Tfive & phi2)
			 | (OP==`SBC_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`SBC_aby & T==`Tfour & phi2)
			 | (OP==`SBC_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`SBC_abx & T==`Tfour & phi2)
			 | (OP==`INC_abx & T==`Tfour & phi2)
			 | (OP==`INC_abx & T==`Tfive & phi1)
			;

assign control[`SB_DB] = (OP==`BRK & T==`Tone & phi2)
			 | (OP==`BRK & T==`Ttwo & phi1)
			 | (OP==`ORA_izx & T==`Tone & phi2)
			 | (OP==`ORA_izx & T==`Ttwo & phi1)
			 | (OP==`ORA_zp & T==`Tone & phi2)
			 | (OP==`ORA_zp & T==`Ttwo & phi1)
			 | (OP==`ASL_zp & T==`Tzero & phi1)
			 | (OP==`ASL_zp & T==`Tone & phi2)
			 | (OP==`ASL_zp & T==`Ttwo & phi1)
			 | (OP==`ASL_zp & T==`Tthree & phi2)
			 | (OP==`ASL_zp & T==`Tfour & phi1)
			 | (OP==`ASL_zp & T==`Tfour & phi2)
			 | (OP==`PHP & T==`Tone & phi2)
			 | (OP==`PHP & T==`Ttwo & phi1)
			 | (OP==`ORA_imm & T==`Tone & phi2)
			 | (OP==`ORA_imm & T==`Ttwo & phi1)
			 | (OP==`ASL & T==`Tone & phi1)
			 | (OP==`ASL & T==`Tone & phi2)
			 | (OP==`ASL & T==`Ttwo & phi1)
			 | (OP==`ASL & T==`Ttwo & phi2)
			 | (OP==`ORA_abs & T==`Tone & phi2)
			 | (OP==`ORA_abs & T==`Ttwo & phi1)
			 | (OP==`ASL_abs & T==`Tzero & phi1)
			 | (OP==`ASL_abs & T==`Tone & phi2)
			 | (OP==`ASL_abs & T==`Ttwo & phi1)
			 | (OP==`ASL_abs & T==`Tfour & phi2)
			 | (OP==`ASL_abs & T==`Tfive & phi1)
			 | (OP==`ASL_abs & T==`Tfive & phi2)
			 | (OP==`BPL_rel & T==`Ttwo & phi1)
			 | (OP==`BPL_rel & T==`Ttwo & phi2)
			 | (OP==`BPL_rel & T==`Tthree & phi1)
			 | (OP==`BPL_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BPL_rel & T==`T1BranchCross & phi2)
			 | (OP==`BPL_rel & T==`T1NoBranch & phi1)
			 | (OP==`BPL_rel & T==`T1NoBranch & phi2)
			 | (OP==`ORA_izy & T==`Tone & phi2)
			 | (OP==`ORA_izy & T==`Ttwo & phi1)
			 | (OP==`ORA_zpx & T==`Tone & phi2)
			 | (OP==`ORA_zpx & T==`Ttwo & phi1)
			 | (OP==`ASL_zpx & T==`Tzero & phi1)
			 | (OP==`ASL_zpx & T==`Tone & phi2)
			 | (OP==`ASL_zpx & T==`Ttwo & phi1)
			 | (OP==`ASL_zpx & T==`Tfour & phi2)
			 | (OP==`ASL_zpx & T==`Tfive & phi1)
			 | (OP==`ASL_zpx & T==`Tfive & phi2)
			 | (OP==`CLC & T==`Tone & phi2)
			 | (OP==`CLC & T==`Ttwo & phi1)
			 | (OP==`ORA_aby & T==`Tone & phi2)
			 | (OP==`ORA_aby & T==`Ttwo & phi1)
			 | (OP==`ORA_abx & T==`Tone & phi2)
			 | (OP==`ORA_abx & T==`Ttwo & phi1)
			 | (OP==`ASL_abx & T==`Tzero & phi1)
			 | (OP==`ASL_abx & T==`Tone & phi2)
			 | (OP==`ASL_abx & T==`Ttwo & phi1)
			 | (OP==`ASL_abx & T==`Tfive & phi2)
			 | (OP==`ASL_abx & T==`Tsix & phi1)
			 | (OP==`ASL_abx & T==`Tsix & phi2)
			 | (OP==`JSR_abs & T==`Tone & phi2)
			 | (OP==`JSR_abs & T==`Ttwo & phi1)
			 | (OP==`JSR_abs & T==`Ttwo & phi2)
			 | (OP==`JSR_abs & T==`Tthree & phi1)
			 | (OP==`AND_izx & T==`Tone & phi2)
			 | (OP==`AND_izx & T==`Ttwo & phi1)
			 | (OP==`BIT_zp & T==`Tone & phi2)
			 | (OP==`BIT_zp & T==`Ttwo & phi1)
			 | (OP==`AND_zp & T==`Tone & phi2)
			 | (OP==`AND_zp & T==`Ttwo & phi1)
			 | (OP==`ROL_zp & T==`Tzero & phi1)
			 | (OP==`ROL_zp & T==`Tone & phi2)
			 | (OP==`ROL_zp & T==`Ttwo & phi1)
			 | (OP==`ROL_zp & T==`Tthree & phi2)
			 | (OP==`ROL_zp & T==`Tfour & phi1)
			 | (OP==`ROL_zp & T==`Tfour & phi2)
			 | (OP==`PLP & T==`Tone & phi2)
			 | (OP==`PLP & T==`Ttwo & phi1)
			 | (OP==`AND_imm & T==`Tone & phi2)
			 | (OP==`AND_imm & T==`Ttwo & phi1)
			 | (OP==`ROL & T==`Tone & phi1)
			 | (OP==`ROL & T==`Tone & phi2)
			 | (OP==`ROL & T==`Ttwo & phi1)
			 | (OP==`ROL & T==`Ttwo & phi2)
			 | (OP==`BIT_abs & T==`Tone & phi2)
			 | (OP==`BIT_abs & T==`Ttwo & phi1)
			 | (OP==`AND_abs & T==`Tone & phi2)
			 | (OP==`AND_abs & T==`Ttwo & phi1)
			 | (OP==`ROL_abs & T==`Tzero & phi1)
			 | (OP==`ROL_abs & T==`Tone & phi2)
			 | (OP==`ROL_abs & T==`Ttwo & phi1)
			 | (OP==`ROL_abs & T==`Tfour & phi2)
			 | (OP==`ROL_abs & T==`Tfive & phi1)
			 | (OP==`ROL_abs & T==`Tfive & phi2)
			 | (OP==`BMI_rel & T==`Ttwo & phi1)
			 | (OP==`BMI_rel & T==`Ttwo & phi2)
			 | (OP==`BMI_rel & T==`Tthree & phi1)
			 | (OP==`BMI_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BMI_rel & T==`T1BranchCross & phi2)
			 | (OP==`BMI_rel & T==`T1NoBranch & phi1)
			 | (OP==`BMI_rel & T==`T1NoBranch & phi2)
			 | (OP==`AND_izy & T==`Tone & phi2)
			 | (OP==`AND_izy & T==`Ttwo & phi1)
			 | (OP==`AND_zpx & T==`Tone & phi2)
			 | (OP==`AND_zpx & T==`Ttwo & phi1)
			 | (OP==`ROL_zpx & T==`Tzero & phi1)
			 | (OP==`ROL_zpx & T==`Tone & phi2)
			 | (OP==`ROL_zpx & T==`Ttwo & phi1)
			 | (OP==`ROL_zpx & T==`Tfour & phi2)
			 | (OP==`ROL_zpx & T==`Tfive & phi1)
			 | (OP==`ROL_zpx & T==`Tfive & phi2)
			 | (OP==`SEC & T==`Tone & phi2)
			 | (OP==`SEC & T==`Ttwo & phi1)
			 | (OP==`AND_aby & T==`Tone & phi2)
			 | (OP==`AND_aby & T==`Ttwo & phi1)
			 | (OP==`AND_abx & T==`Tone & phi2)
			 | (OP==`AND_abx & T==`Ttwo & phi1)
			 | (OP==`ROL_abx & T==`Tzero & phi1)
			 | (OP==`ROL_abx & T==`Tone & phi2)
			 | (OP==`ROL_abx & T==`Ttwo & phi1)
			 | (OP==`ROL_abx & T==`Tfive & phi2)
			 | (OP==`ROL_abx & T==`Tsix & phi1)
			 | (OP==`ROL_abx & T==`Tsix & phi2)
			 | (OP==`RTI & T==`Tone & phi2)
			 | (OP==`RTI & T==`Ttwo & phi1)
			 | (OP==`EOR_izx & T==`Tone & phi2)
			 | (OP==`EOR_izx & T==`Ttwo & phi1)
			 | (OP==`EOR_zp & T==`Tone & phi2)
			 | (OP==`EOR_zp & T==`Ttwo & phi1)
			 | (OP==`LSR_zp & T==`Tzero & phi1)
			 | (OP==`LSR_zp & T==`Tone & phi2)
			 | (OP==`LSR_zp & T==`Ttwo & phi1)
			 | (OP==`LSR_zp & T==`Tfour & phi2)
			 | (OP==`PHA & T==`Tone & phi2)
			 | (OP==`PHA & T==`Ttwo & phi1)
			 | (OP==`EOR_imm & T==`Tone & phi2)
			 | (OP==`EOR_imm & T==`Ttwo & phi1)
			 | (OP==`LSR & T==`Tone & phi1)
			 | (OP==`LSR & T==`Tone & phi2)
			 | (OP==`LSR & T==`Ttwo & phi1)
			 | (OP==`LSR & T==`Ttwo & phi2)
			 | (OP==`JMP_abs & T==`Tone & phi2)
			 | (OP==`JMP_abs & T==`Ttwo & phi1)
			 | (OP==`EOR_abs & T==`Tone & phi2)
			 | (OP==`EOR_abs & T==`Ttwo & phi1)
			 | (OP==`LSR_abs & T==`Tzero & phi1)
			 | (OP==`LSR_abs & T==`Tone & phi2)
			 | (OP==`LSR_abs & T==`Ttwo & phi1)
			 | (OP==`LSR_abs & T==`Tfive & phi2)
			 | (OP==`BVC_rel & T==`Ttwo & phi1)
			 | (OP==`BVC_rel & T==`Ttwo & phi2)
			 | (OP==`BVC_rel & T==`Tthree & phi1)
			 | (OP==`BVC_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BVC_rel & T==`T1BranchCross & phi2)
			 | (OP==`BVC_rel & T==`T1NoBranch & phi1)
			 | (OP==`BVC_rel & T==`T1NoBranch & phi2)
			 | (OP==`EOR_izy & T==`Tone & phi2)
			 | (OP==`EOR_izy & T==`Ttwo & phi1)
			 | (OP==`EOR_zpx & T==`Tone & phi2)
			 | (OP==`EOR_zpx & T==`Ttwo & phi1)
			 | (OP==`LSR_zpx & T==`Tzero & phi1)
			 | (OP==`LSR_zpx & T==`Tone & phi2)
			 | (OP==`LSR_zpx & T==`Ttwo & phi1)
			 | (OP==`LSR_zpx & T==`Tfive & phi2)
			 | (OP==`CLI & T==`Tone & phi2)
			 | (OP==`CLI & T==`Ttwo & phi1)
			 | (OP==`EOR_aby & T==`Tone & phi2)
			 | (OP==`EOR_aby & T==`Ttwo & phi1)
			 | (OP==`EOR_abx & T==`Tone & phi2)
			 | (OP==`EOR_abx & T==`Ttwo & phi1)
			 | (OP==`LSR_abx & T==`Tzero & phi1)
			 | (OP==`LSR_abx & T==`Tone & phi2)
			 | (OP==`LSR_abx & T==`Ttwo & phi1)
			 | (OP==`LSR_abx & T==`Tsix & phi2)
			 | (OP==`RTS & T==`Tone & phi2)
			 | (OP==`RTS & T==`Ttwo & phi1)
			 | (OP==`ADC_izx & T==`Tone & phi2)
			 | (OP==`ADC_izx & T==`Ttwo & phi1)
			 | (OP==`ADC_zp & T==`Tone & phi2)
			 | (OP==`ADC_zp & T==`Ttwo & phi1)
			 | (OP==`ROR_zp & T==`Tzero & phi1)
			 | (OP==`ROR_zp & T==`Tone & phi2)
			 | (OP==`ROR_zp & T==`Ttwo & phi1)
			 | (OP==`ROR_zp & T==`Tfour & phi2)
			 | (OP==`PLA & T==`Tzero & phi2)
			 | (OP==`PLA & T==`Tone & phi1)
			 | (OP==`PLA & T==`Tone & phi2)
			 | (OP==`PLA & T==`Ttwo & phi1)
			 | (OP==`ADC_imm & T==`Tone & phi2)
			 | (OP==`ADC_imm & T==`Ttwo & phi1)
			 | (OP==`ROR & T==`Tone & phi1)
			 | (OP==`ROR & T==`Tone & phi2)
			 | (OP==`ROR & T==`Ttwo & phi1)
			 | (OP==`ROR & T==`Ttwo & phi2)
			 | (OP==`JMP_zp & T==`Tone & phi2)
			 | (OP==`JMP_zp & T==`Ttwo & phi1)
			 | (OP==`ADC_abs & T==`Tone & phi2)
			 | (OP==`ADC_abs & T==`Ttwo & phi1)
			 | (OP==`ROR_abs & T==`Tzero & phi1)
			 | (OP==`ROR_abs & T==`Tone & phi2)
			 | (OP==`ROR_abs & T==`Ttwo & phi1)
			 | (OP==`ROR_abs & T==`Tfive & phi2)
			 | (OP==`BVS_rel & T==`Ttwo & phi1)
			 | (OP==`BVS_rel & T==`Ttwo & phi2)
			 | (OP==`BVS_rel & T==`Tthree & phi1)
			 | (OP==`BVS_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BVS_rel & T==`T1BranchCross & phi2)
			 | (OP==`BVS_rel & T==`T1NoBranch & phi1)
			 | (OP==`BVS_rel & T==`T1NoBranch & phi2)
			 | (OP==`ADC_izy & T==`Tone & phi2)
			 | (OP==`ADC_izy & T==`Ttwo & phi1)
			 | (OP==`ADC_zpx & T==`Tone & phi2)
			 | (OP==`ADC_zpx & T==`Ttwo & phi1)
			 | (OP==`ROR_zpx & T==`Tzero & phi1)
			 | (OP==`ROR_zpx & T==`Tone & phi2)
			 | (OP==`ROR_zpx & T==`Ttwo & phi1)
			 | (OP==`ROR_zpx & T==`Tfive & phi2)
			 | (OP==`SEI & T==`Tone & phi2)
			 | (OP==`SEI & T==`Ttwo & phi1)
			 | (OP==`ADC_aby & T==`Tone & phi2)
			 | (OP==`ADC_aby & T==`Ttwo & phi1)
			 | (OP==`ADC_abx & T==`Tone & phi2)
			 | (OP==`ADC_abx & T==`Ttwo & phi1)
			 | (OP==`ROR_abx & T==`Tzero & phi1)
			 | (OP==`ROR_abx & T==`Tone & phi2)
			 | (OP==`ROR_abx & T==`Ttwo & phi1)
			 | (OP==`ROR_abx & T==`Tsix & phi2)
			 | (OP==`STA_izx & T==`Tone & phi2)
			 | (OP==`STA_izx & T==`Ttwo & phi1)
			 | (OP==`STY_zp & T==`Tzero & phi1)
			 | (OP==`STY_zp & T==`Tone & phi2)
			 | (OP==`STY_zp & T==`Ttwo & phi1)
			 | (OP==`STY_zp & T==`Ttwo & phi2)
			 | (OP==`STA_zp & T==`Tone & phi2)
			 | (OP==`STA_zp & T==`Ttwo & phi1)
			 | (OP==`STX_zp & T==`Tzero & phi1)
			 | (OP==`STX_zp & T==`Tone & phi2)
			 | (OP==`STX_zp & T==`Ttwo & phi1)
			 | (OP==`STX_zp & T==`Ttwo & phi2)
			 | (OP==`DEY & T==`Tone & phi2)
			 | (OP==`DEY & T==`Ttwo & phi1)
			 | (OP==`TXA & T==`Tone & phi1)
			 | (OP==`TXA & T==`Tone & phi2)
			 | (OP==`TXA & T==`Ttwo & phi1)
			 | (OP==`TXA & T==`Ttwo & phi2)
			 | (OP==`STY_abs & T==`Tzero & phi1)
			 | (OP==`STY_abs & T==`Tone & phi2)
			 | (OP==`STY_abs & T==`Ttwo & phi1)
			 | (OP==`STY_abs & T==`Tthree & phi2)
			 | (OP==`STA_abs & T==`Tone & phi2)
			 | (OP==`STA_abs & T==`Ttwo & phi1)
			 | (OP==`STX_abs & T==`Tzero & phi1)
			 | (OP==`STX_abs & T==`Tone & phi2)
			 | (OP==`STX_abs & T==`Ttwo & phi1)
			 | (OP==`STX_abs & T==`Tthree & phi2)
			 | (OP==`BCC_rel & T==`Ttwo & phi1)
			 | (OP==`BCC_rel & T==`Ttwo & phi2)
			 | (OP==`BCC_rel & T==`Tthree & phi1)
			 | (OP==`BCC_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BCC_rel & T==`T1BranchCross & phi2)
			 | (OP==`BCC_rel & T==`T1NoBranch & phi1)
			 | (OP==`BCC_rel & T==`T1NoBranch & phi2)
			 | (OP==`STA_izy & T==`Tone & phi2)
			 | (OP==`STA_izy & T==`Ttwo & phi1)
			 | (OP==`STY_zpx & T==`Tzero & phi1)
			 | (OP==`STY_zpx & T==`Tone & phi2)
			 | (OP==`STY_zpx & T==`Ttwo & phi1)
			 | (OP==`STY_zpx & T==`Tthree & phi2)
			 | (OP==`STA_zpx & T==`Tone & phi2)
			 | (OP==`STA_zpx & T==`Ttwo & phi1)
			 | (OP==`STX_zpy & T==`Tzero & phi1)
			 | (OP==`STX_zpy & T==`Tone & phi2)
			 | (OP==`STX_zpy & T==`Ttwo & phi1)
			 | (OP==`STX_zpy & T==`Tthree & phi2)
			 | (OP==`TYA & T==`Tone & phi1)
			 | (OP==`TYA & T==`Tone & phi2)
			 | (OP==`TYA & T==`Ttwo & phi1)
			 | (OP==`TYA & T==`Ttwo & phi2)
			 | (OP==`STA_aby & T==`Tone & phi2)
			 | (OP==`STA_aby & T==`Ttwo & phi1)
			 | (OP==`TXS & T==`Tone & phi1)
			 | (OP==`TXS & T==`Tone & phi2)
			 | (OP==`TXS & T==`Ttwo & phi1)
			 | (OP==`STA_abx & T==`Tone & phi2)
			 | (OP==`STA_abx & T==`Ttwo & phi1)
			 | (OP==`LDY_imm & T==`Tone & phi1)
			 | (OP==`LDY_imm & T==`Tone & phi2)
			 | (OP==`LDY_imm & T==`Ttwo & phi1)
			 | (OP==`LDY_imm & T==`Ttwo & phi2)
			 | (OP==`LDA_izx & T==`Tzero & phi2)
			 | (OP==`LDA_izx & T==`Tone & phi1)
			 | (OP==`LDA_izx & T==`Tone & phi2)
			 | (OP==`LDA_izx & T==`Ttwo & phi1)
			 | (OP==`LDX_imm & T==`Tone & phi1)
			 | (OP==`LDX_imm & T==`Tone & phi2)
			 | (OP==`LDX_imm & T==`Ttwo & phi1)
			 | (OP==`LDX_imm & T==`Ttwo & phi2)
			 | (OP==`LDY_zp & T==`Tzero & phi2)
			 | (OP==`LDY_zp & T==`Tone & phi1)
			 | (OP==`LDY_zp & T==`Tone & phi2)
			 | (OP==`LDY_zp & T==`Ttwo & phi1)
			 | (OP==`LDA_zp & T==`Tzero & phi2)
			 | (OP==`LDA_zp & T==`Tone & phi1)
			 | (OP==`LDA_zp & T==`Tone & phi2)
			 | (OP==`LDA_zp & T==`Ttwo & phi1)
			 | (OP==`LDX_zp & T==`Tzero & phi2)
			 | (OP==`LDX_zp & T==`Tone & phi1)
			 | (OP==`LDX_zp & T==`Tone & phi2)
			 | (OP==`LDX_zp & T==`Ttwo & phi1)
			 | (OP==`TAY & T==`Tone & phi1)
			 | (OP==`TAY & T==`Tone & phi2)
			 | (OP==`TAY & T==`Ttwo & phi1)
			 | (OP==`TAY & T==`Ttwo & phi2)
			 | (OP==`LDA_imm & T==`Tone & phi1)
			 | (OP==`LDA_imm & T==`Tone & phi2)
			 | (OP==`LDA_imm & T==`Ttwo & phi1)
			 | (OP==`LDA_imm & T==`Ttwo & phi2)
			 | (OP==`TAX & T==`Tone & phi1)
			 | (OP==`TAX & T==`Tone & phi2)
			 | (OP==`TAX & T==`Ttwo & phi1)
			 | (OP==`TAX & T==`Ttwo & phi2)
			 | (OP==`LDY_abs & T==`Tzero & phi2)
			 | (OP==`LDY_abs & T==`Tone & phi1)
			 | (OP==`LDY_abs & T==`Tone & phi2)
			 | (OP==`LDY_abs & T==`Ttwo & phi1)
			 | (OP==`LDA_abs & T==`Tzero & phi2)
			 | (OP==`LDA_abs & T==`Tone & phi1)
			 | (OP==`LDA_abs & T==`Tone & phi2)
			 | (OP==`LDA_abs & T==`Ttwo & phi1)
			 | (OP==`LDX_abs & T==`Tzero & phi2)
			 | (OP==`LDX_abs & T==`Tone & phi1)
			 | (OP==`LDX_abs & T==`Tone & phi2)
			 | (OP==`LDX_abs & T==`Ttwo & phi1)
			 | (OP==`BCS_rel & T==`Ttwo & phi1)
			 | (OP==`BCS_rel & T==`Ttwo & phi2)
			 | (OP==`BCS_rel & T==`Tthree & phi1)
			 | (OP==`BCS_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BCS_rel & T==`T1BranchCross & phi2)
			 | (OP==`BCS_rel & T==`T1NoBranch & phi1)
			 | (OP==`BCS_rel & T==`T1NoBranch & phi2)
			 | (OP==`LDA_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`LDA_izy & T==`TzeroCrossPg & phi2)
			 | (OP==`LDA_izy & T==`Tone & phi1)
			 | (OP==`LDA_izy & T==`Tone & phi2)
			 | (OP==`LDA_izy & T==`Ttwo & phi1)
			 | (OP==`LDY_zpx & T==`Tzero & phi2)
			 | (OP==`LDY_zpx & T==`Tone & phi1)
			 | (OP==`LDY_zpx & T==`Tone & phi2)
			 | (OP==`LDY_zpx & T==`Ttwo & phi1)
			 | (OP==`LDA_zpx & T==`Tzero & phi2)
			 | (OP==`LDA_zpx & T==`Tone & phi1)
			 | (OP==`LDA_zpx & T==`Tone & phi2)
			 | (OP==`LDA_zpx & T==`Ttwo & phi1)
			 | (OP==`LDX_zpy & T==`Tzero & phi2)
			 | (OP==`LDX_zpy & T==`Tone & phi1)
			 | (OP==`LDX_zpy & T==`Tone & phi2)
			 | (OP==`LDX_zpy & T==`Ttwo & phi1)
			 | (OP==`CLV & T==`Tone & phi2)
			 | (OP==`CLV & T==`Ttwo & phi1)
			 | (OP==`LDA_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`LDA_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`LDA_aby & T==`Tone & phi1)
			 | (OP==`LDA_aby & T==`Tone & phi2)
			 | (OP==`LDA_aby & T==`Ttwo & phi1)
			 | (OP==`TSX & T==`Tone & phi1)
			 | (OP==`TSX & T==`Tone & phi2)
			 | (OP==`TSX & T==`Ttwo & phi1)
			 | (OP==`TSX & T==`Ttwo & phi2)
			 | (OP==`LDY_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`LDY_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`LDY_abx & T==`Tone & phi1)
			 | (OP==`LDY_abx & T==`Tone & phi2)
			 | (OP==`LDY_abx & T==`Ttwo & phi1)
			 | (OP==`LDA_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`LDA_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`LDA_abx & T==`Tone & phi1)
			 | (OP==`LDA_abx & T==`Tone & phi2)
			 | (OP==`LDA_abx & T==`Ttwo & phi1)
			 | (OP==`LDX_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`LDX_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`LDX_aby & T==`Tone & phi1)
			 | (OP==`LDX_aby & T==`Tone & phi2)
			 | (OP==`LDX_aby & T==`Ttwo & phi1)
			 | (OP==`CPY_imm & T==`Tone & phi2)
			 | (OP==`CPY_imm & T==`Ttwo & phi1)
			 | (OP==`CMP_izx & T==`Tone & phi2)
			 | (OP==`CMP_izx & T==`Ttwo & phi1)
			 | (OP==`CPY_zp & T==`Tone & phi2)
			 | (OP==`CPY_zp & T==`Ttwo & phi1)
			 | (OP==`CMP_zp & T==`Tone & phi2)
			 | (OP==`CMP_zp & T==`Ttwo & phi1)
			 | (OP==`DEC_zp & T==`Tzero & phi1)
			 | (OP==`DEC_zp & T==`Tone & phi2)
			 | (OP==`DEC_zp & T==`Ttwo & phi1)
			 | (OP==`DEC_zp & T==`Tfour & phi2)
			 | (OP==`INY & T==`Tone & phi2)
			 | (OP==`INY & T==`Ttwo & phi1)
			 | (OP==`CMP_imm & T==`Tone & phi2)
			 | (OP==`CMP_imm & T==`Ttwo & phi1)
			 | (OP==`DEX & T==`Tone & phi2)
			 | (OP==`DEX & T==`Ttwo & phi1)
			 | (OP==`CPY_abs & T==`Tone & phi2)
			 | (OP==`CPY_abs & T==`Ttwo & phi1)
			 | (OP==`CMP_abs & T==`Tone & phi2)
			 | (OP==`CMP_abs & T==`Ttwo & phi1)
			 | (OP==`DEC_abs & T==`Tzero & phi1)
			 | (OP==`DEC_abs & T==`Tone & phi2)
			 | (OP==`DEC_abs & T==`Ttwo & phi1)
			 | (OP==`DEC_abs & T==`Tfive & phi2)
			 | (OP==`BNE_rel & T==`Ttwo & phi1)
			 | (OP==`BNE_rel & T==`Ttwo & phi2)
			 | (OP==`BNE_rel & T==`Tthree & phi1)
			 | (OP==`BNE_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BNE_rel & T==`T1BranchCross & phi2)
			 | (OP==`BNE_rel & T==`T1NoBranch & phi1)
			 | (OP==`BNE_rel & T==`T1NoBranch & phi2)
			 | (OP==`CMP_izy & T==`Tone & phi2)
			 | (OP==`CMP_izy & T==`Ttwo & phi1)
			 | (OP==`CMP_zpx & T==`Tone & phi2)
			 | (OP==`CMP_zpx & T==`Ttwo & phi1)
			 | (OP==`DEC_zpx & T==`Tzero & phi1)
			 | (OP==`DEC_zpx & T==`Tone & phi2)
			 | (OP==`DEC_zpx & T==`Ttwo & phi1)
			 | (OP==`DEC_zpx & T==`Tfive & phi2)
			 | (OP==`CLD & T==`Tone & phi2)
			 | (OP==`CLD & T==`Ttwo & phi1)
			 | (OP==`CMP_aby & T==`Tone & phi2)
			 | (OP==`CMP_aby & T==`Ttwo & phi1)
			 | (OP==`CMP_abx & T==`Tone & phi2)
			 | (OP==`CMP_abx & T==`Ttwo & phi1)
			 | (OP==`DEC_abx & T==`Tzero & phi1)
			 | (OP==`DEC_abx & T==`Tone & phi2)
			 | (OP==`DEC_abx & T==`Ttwo & phi1)
			 | (OP==`DEC_abx & T==`Tsix & phi2)
			 | (OP==`CPX_imm & T==`Tone & phi2)
			 | (OP==`CPX_imm & T==`Ttwo & phi1)
			 | (OP==`SBC_izx & T==`Tone & phi2)
			 | (OP==`SBC_izx & T==`Ttwo & phi1)
			 | (OP==`CPX_zp & T==`Tone & phi2)
			 | (OP==`CPX_zp & T==`Ttwo & phi1)
			 | (OP==`SBC_zp & T==`Tone & phi2)
			 | (OP==`SBC_zp & T==`Ttwo & phi1)
			 | (OP==`INC_zp & T==`Tzero & phi1)
			 | (OP==`INC_zp & T==`Tone & phi2)
			 | (OP==`INC_zp & T==`Ttwo & phi1)
			 | (OP==`INC_zp & T==`Tfour & phi2)
			 | (OP==`INX & T==`Tone & phi2)
			 | (OP==`INX & T==`Ttwo & phi1)
			 | (OP==`SBC_imm & T==`Tone & phi2)
			 | (OP==`SBC_imm & T==`Ttwo & phi1)
			 | (OP==`NOP & T==`Tone & phi2)
			 | (OP==`NOP & T==`Ttwo & phi1)
			 | (OP==`CPX_abs & T==`Tone & phi2)
			 | (OP==`CPX_abs & T==`Ttwo & phi1)
			 | (OP==`SBC_abs & T==`Tone & phi2)
			 | (OP==`SBC_abs & T==`Ttwo & phi1)
			 | (OP==`INC_abs & T==`Tzero & phi1)
			 | (OP==`INC_abs & T==`Tone & phi2)
			 | (OP==`INC_abs & T==`Ttwo & phi1)
			 | (OP==`INC_abs & T==`Tfive & phi2)
			 | (OP==`BEQ_rel & T==`Ttwo & phi1)
			 | (OP==`BEQ_rel & T==`Ttwo & phi2)
			 | (OP==`BEQ_rel & T==`Tthree & phi1)
			 | (OP==`BEQ_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BEQ_rel & T==`T1BranchCross & phi2)
			 | (OP==`BEQ_rel & T==`T1NoBranch & phi1)
			 | (OP==`BEQ_rel & T==`T1NoBranch & phi2)
			 | (OP==`SBC_izy & T==`Tone & phi2)
			 | (OP==`SBC_izy & T==`Ttwo & phi1)
			 | (OP==`SBC_zpx & T==`Tone & phi2)
			 | (OP==`SBC_zpx & T==`Ttwo & phi1)
			 | (OP==`INC_zpx & T==`Tzero & phi1)
			 | (OP==`INC_zpx & T==`Tone & phi2)
			 | (OP==`INC_zpx & T==`Ttwo & phi1)
			 | (OP==`INC_zpx & T==`Tfive & phi2)
			 | (OP==`SED & T==`Tone & phi2)
			 | (OP==`SED & T==`Ttwo & phi1)
			 | (OP==`SBC_aby & T==`Tone & phi2)
			 | (OP==`SBC_aby & T==`Ttwo & phi1)
			 | (OP==`SBC_abx & T==`Tone & phi2)
			 | (OP==`SBC_abx & T==`Ttwo & phi1)
			 | (OP==`INC_abx & T==`Tzero & phi1)
			 | (OP==`INC_abx & T==`Tone & phi2)
			 | (OP==`INC_abx & T==`Ttwo & phi1)
			 | (OP==`INC_abx & T==`Tsix & phi2)
			;

assign control[`O_ADL0] = (OP==`BRK & (activeInt == `RST_i | activeInt == `IRQ_i | activeInt == `NMI_i | activeInt == `NONE) &
			((T==`Tfive & phi2) | (T==`Tsix & phi1)));

assign control[`O_ADL1] = (OP==`BRK & activeInt == `RST_i & ((T==`Tfive & phi2) |
			(T==`Tsix) |
			(T==`Tzero& phi1)));

assign control[`O_ADL2] = (OP==`BRK & activeInt == `NMI_i & ((T==`Tfive & phi2) |
			(T==`Tsix) |
			(T==`Tzero & phi1)));

assign control[`S_ADL] = (OP==`BRK & T==`Ttwo & phi2)
			 | (OP==`BRK & T==`Tthree & phi1)
			 | (OP==`PHP & T==`Tzero & phi1)
			 | (OP==`PHP & T==`Ttwo & phi2)
			 | (OP==`JSR_abs & T==`Tzero & phi2)
			 | (OP==`JSR_abs & T==`Tone & phi1)
			 | (OP==`JSR_abs & T==`Ttwo & phi2)
			 | (OP==`JSR_abs & T==`Tthree & phi1)
			 | (OP==`PLP & T==`Ttwo & phi2)
			 | (OP==`PLP & T==`Tthree & phi1)
			 | (OP==`RTI & T==`Ttwo & phi2)
			 | (OP==`RTI & T==`Tthree & phi1)
			 | (OP==`PHA & T==`Tzero & phi1)
			 | (OP==`PHA & T==`Ttwo & phi2)
			 | (OP==`RTS & T==`Ttwo & phi2)
			 | (OP==`RTS & T==`Tthree & phi1)
			 | (OP==`PLA & T==`Ttwo & phi2)
			 | (OP==`PLA & T==`Tthree & phi1)
			;

assign control[`SB_S] = (OP==`BRK & T==`Tsix & phi1)
			 | (OP==`PHP & T==`Tone & phi1)
			 | (OP==`JSR_abs & T==`Tone & phi1)
			 | (OP==`JSR_abs & T==`Tthree & phi1)
			 | (OP==`PLP & T==`Tzero & phi1)
			 | (OP==`RTI & T==`Tzero & phi1)
			 | (OP==`PHA & T==`Tone & phi1)
			 | (OP==`RTS & T==`Tfive & phi1)
			 | (OP==`PLA & T==`Tzero & phi1)
			 | (OP==`TXS & T==`Tone & phi1)
			;

assign control[`S_S] = (OP==`BRK & T==`Tzero & phi1)
			 | (OP==`BRK & T==`Tone & phi1)
			 | (OP==`BRK & T==`Ttwo & phi1)
			 | (OP==`BRK & T==`Tthree & phi1)
			 | (OP==`BRK & T==`Tfour & phi1)
			 | (OP==`BRK & T==`Tfive & phi1)
			 | (OP==`ORA_izx & T==`Tzero & phi1)
			 | (OP==`ORA_izx & T==`Tone & phi1)
			 | (OP==`ORA_izx & T==`Ttwo & phi1)
			 | (OP==`ORA_izx & T==`Tthree & phi1)
			 | (OP==`ORA_izx & T==`Tfour & phi1)
			 | (OP==`ORA_izx & T==`Tfive & phi1)
			 | (OP==`ORA_zp & T==`Tzero & phi1)
			 | (OP==`ORA_zp & T==`Tone & phi1)
			 | (OP==`ORA_zp & T==`Ttwo & phi1)
			 | (OP==`ASL_zp & T==`Tzero & phi1)
			 | (OP==`ASL_zp & T==`Tone & phi1)
			 | (OP==`ASL_zp & T==`Ttwo & phi1)
			 | (OP==`ASL_zp & T==`Tthree & phi1)
			 | (OP==`ASL_zp & T==`Tfour & phi1)
			 | (OP==`PHP & T==`Tzero & phi1)
			 | (OP==`PHP & T==`Ttwo & phi1)
			 | (OP==`ORA_imm & T==`Tone & phi1)
			 | (OP==`ORA_imm & T==`Ttwo & phi1)
			 | (OP==`ASL & T==`Tone & phi1)
			 | (OP==`ASL & T==`Ttwo & phi1)
			 | (OP==`ORA_abs & T==`Tzero & phi1)
			 | (OP==`ORA_abs & T==`Tone & phi1)
			 | (OP==`ORA_abs & T==`Ttwo & phi1)
			 | (OP==`ORA_abs & T==`Tthree & phi1)
			 | (OP==`ASL_abs & T==`Tzero & phi1)
			 | (OP==`ASL_abs & T==`Tone & phi1)
			 | (OP==`ASL_abs & T==`Ttwo & phi1)
			 | (OP==`ASL_abs & T==`Tthree & phi1)
			 | (OP==`ASL_abs & T==`Tfour & phi1)
			 | (OP==`ASL_abs & T==`Tfive & phi1)
			 | (OP==`BPL_rel & T==`Tzero & phi1)
			 | (OP==`BPL_rel & T==`Ttwo & phi1)
			 | (OP==`BPL_rel & T==`Tthree & phi1)
			 | (OP==`BPL_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BPL_rel & T==`T1BranchCross & phi1)
			 | (OP==`BPL_rel & T==`T1NoBranch & phi1)
			 | (OP==`ORA_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`ORA_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ORA_izy & T==`Tone & phi1)
			 | (OP==`ORA_izy & T==`Ttwo & phi1)
			 | (OP==`ORA_izy & T==`Tthree & phi1)
			 | (OP==`ORA_izy & T==`Tfour & phi1)
			 | (OP==`ORA_izy & T==`Tfive & phi1)
			 | (OP==`ORA_zpx & T==`Tzero & phi1)
			 | (OP==`ORA_zpx & T==`Tone & phi1)
			 | (OP==`ORA_zpx & T==`Ttwo & phi1)
			 | (OP==`ORA_zpx & T==`Tthree & phi1)
			 | (OP==`ASL_zpx & T==`Tzero & phi1)
			 | (OP==`ASL_zpx & T==`Tone & phi1)
			 | (OP==`ASL_zpx & T==`Ttwo & phi1)
			 | (OP==`ASL_zpx & T==`Tthree & phi1)
			 | (OP==`ASL_zpx & T==`Tfour & phi1)
			 | (OP==`ASL_zpx & T==`Tfive & phi1)
			 | (OP==`CLC & T==`Tone & phi1)
			 | (OP==`CLC & T==`Ttwo & phi1)
			 | (OP==`ORA_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ORA_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`ORA_aby & T==`Tone & phi1)
			 | (OP==`ORA_aby & T==`Ttwo & phi1)
			 | (OP==`ORA_aby & T==`Tthree & phi1)
			 | (OP==`ORA_aby & T==`Tfour & phi1)
			 | (OP==`ORA_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ORA_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`ORA_abx & T==`Tone & phi1)
			 | (OP==`ORA_abx & T==`Ttwo & phi1)
			 | (OP==`ORA_abx & T==`Tthree & phi1)
			 | (OP==`ORA_abx & T==`Tfour & phi1)
			 | (OP==`ASL_abx & T==`Tzero & phi1)
			 | (OP==`ASL_abx & T==`Tone & phi1)
			 | (OP==`ASL_abx & T==`Ttwo & phi1)
			 | (OP==`ASL_abx & T==`Tthree & phi1)
			 | (OP==`ASL_abx & T==`Tfour & phi1)
			 | (OP==`ASL_abx & T==`Tfive & phi1)
			 | (OP==`ASL_abx & T==`Tsix & phi1)
			 | (OP==`JSR_abs & T==`Tzero & phi1)
			 | (OP==`JSR_abs & T==`Ttwo & phi1)
			 | (OP==`JSR_abs & T==`Tfour & phi1)
			 | (OP==`JSR_abs & T==`Tfive & phi1)
			 | (OP==`AND_izx & T==`Tzero & phi1)
			 | (OP==`AND_izx & T==`Tone & phi1)
			 | (OP==`AND_izx & T==`Ttwo & phi1)
			 | (OP==`AND_izx & T==`Tthree & phi1)
			 | (OP==`AND_izx & T==`Tfour & phi1)
			 | (OP==`AND_izx & T==`Tfive & phi1)
			 | (OP==`BIT_zp & T==`Tzero & phi1)
			 | (OP==`BIT_zp & T==`Tone & phi1)
			 | (OP==`BIT_zp & T==`Ttwo & phi1)
			 | (OP==`AND_zp & T==`Tzero & phi1)
			 | (OP==`AND_zp & T==`Tone & phi1)
			 | (OP==`AND_zp & T==`Ttwo & phi1)
			 | (OP==`ROL_zp & T==`Tzero & phi1)
			 | (OP==`ROL_zp & T==`Tone & phi1)
			 | (OP==`ROL_zp & T==`Ttwo & phi1)
			 | (OP==`ROL_zp & T==`Tthree & phi1)
			 | (OP==`ROL_zp & T==`Tfour & phi1)
			 | (OP==`PLP & T==`Tone & phi1)
			 | (OP==`PLP & T==`Ttwo & phi1)
			 | (OP==`PLP & T==`Tthree & phi1)
			 | (OP==`AND_imm & T==`Tone & phi1)
			 | (OP==`AND_imm & T==`Ttwo & phi1)
			 | (OP==`ROL & T==`Tone & phi1)
			 | (OP==`ROL & T==`Ttwo & phi1)
			 | (OP==`BIT_abs & T==`Tzero & phi1)
			 | (OP==`BIT_abs & T==`Tone & phi1)
			 | (OP==`BIT_abs & T==`Ttwo & phi1)
			 | (OP==`BIT_abs & T==`Tthree & phi1)
			 | (OP==`AND_abs & T==`Tzero & phi1)
			 | (OP==`AND_abs & T==`Tone & phi1)
			 | (OP==`AND_abs & T==`Ttwo & phi1)
			 | (OP==`AND_abs & T==`Tthree & phi1)
			 | (OP==`ROL_abs & T==`Tzero & phi1)
			 | (OP==`ROL_abs & T==`Tone & phi1)
			 | (OP==`ROL_abs & T==`Ttwo & phi1)
			 | (OP==`ROL_abs & T==`Tthree & phi1)
			 | (OP==`ROL_abs & T==`Tfour & phi1)
			 | (OP==`ROL_abs & T==`Tfive & phi1)
			 | (OP==`BMI_rel & T==`Tzero & phi1)
			 | (OP==`BMI_rel & T==`Ttwo & phi1)
			 | (OP==`BMI_rel & T==`Tthree & phi1)
			 | (OP==`BMI_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BMI_rel & T==`T1BranchCross & phi1)
			 | (OP==`BMI_rel & T==`T1NoBranch & phi1)
			 | (OP==`AND_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`AND_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`AND_izy & T==`Tone & phi1)
			 | (OP==`AND_izy & T==`Ttwo & phi1)
			 | (OP==`AND_izy & T==`Tthree & phi1)
			 | (OP==`AND_izy & T==`Tfour & phi1)
			 | (OP==`AND_izy & T==`Tfive & phi1)
			 | (OP==`AND_zpx & T==`Tzero & phi1)
			 | (OP==`AND_zpx & T==`Tone & phi1)
			 | (OP==`AND_zpx & T==`Ttwo & phi1)
			 | (OP==`AND_zpx & T==`Tthree & phi1)
			 | (OP==`ROL_zpx & T==`Tzero & phi1)
			 | (OP==`ROL_zpx & T==`Tone & phi1)
			 | (OP==`ROL_zpx & T==`Ttwo & phi1)
			 | (OP==`ROL_zpx & T==`Tthree & phi1)
			 | (OP==`ROL_zpx & T==`Tfour & phi1)
			 | (OP==`ROL_zpx & T==`Tfive & phi1)
			 | (OP==`SEC & T==`Tone & phi1)
			 | (OP==`SEC & T==`Ttwo & phi1)
			 | (OP==`AND_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`AND_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`AND_aby & T==`Tone & phi1)
			 | (OP==`AND_aby & T==`Ttwo & phi1)
			 | (OP==`AND_aby & T==`Tthree & phi1)
			 | (OP==`AND_aby & T==`Tfour & phi1)
			 | (OP==`AND_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`AND_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`AND_abx & T==`Tone & phi1)
			 | (OP==`AND_abx & T==`Ttwo & phi1)
			 | (OP==`AND_abx & T==`Tthree & phi1)
			 | (OP==`AND_abx & T==`Tfour & phi1)
			 | (OP==`ROL_abx & T==`Tzero & phi1)
			 | (OP==`ROL_abx & T==`Tone & phi1)
			 | (OP==`ROL_abx & T==`Ttwo & phi1)
			 | (OP==`ROL_abx & T==`Tthree & phi1)
			 | (OP==`ROL_abx & T==`Tfour & phi1)
			 | (OP==`ROL_abx & T==`Tfive & phi1)
			 | (OP==`ROL_abx & T==`Tsix & phi1)
			 | (OP==`RTI & T==`Tone & phi1)
			 | (OP==`RTI & T==`Ttwo & phi1)
			 | (OP==`RTI & T==`Tthree & phi1)
			 | (OP==`RTI & T==`Tfour & phi1)
			 | (OP==`RTI & T==`Tfive & phi1)
			 | (OP==`EOR_izx & T==`Tzero & phi1)
			 | (OP==`EOR_izx & T==`Tone & phi1)
			 | (OP==`EOR_izx & T==`Ttwo & phi1)
			 | (OP==`EOR_izx & T==`Tthree & phi1)
			 | (OP==`EOR_izx & T==`Tfour & phi1)
			 | (OP==`EOR_izx & T==`Tfive & phi1)
			 | (OP==`EOR_zp & T==`Tzero & phi1)
			 | (OP==`EOR_zp & T==`Tone & phi1)
			 | (OP==`EOR_zp & T==`Ttwo & phi1)
			 | (OP==`LSR_zp & T==`Tzero & phi1)
			 | (OP==`LSR_zp & T==`Tone & phi1)
			 | (OP==`LSR_zp & T==`Ttwo & phi1)
			 | (OP==`LSR_zp & T==`Tthree & phi1)
			 | (OP==`LSR_zp & T==`Tfour & phi1)
			 | (OP==`PHA & T==`Tzero & phi1)
			 | (OP==`PHA & T==`Ttwo & phi1)
			 | (OP==`EOR_imm & T==`Tone & phi1)
			 | (OP==`EOR_imm & T==`Ttwo & phi1)
			 | (OP==`LSR & T==`Tone & phi1)
			 | (OP==`LSR & T==`Ttwo & phi1)
			 | (OP==`JMP_abs & T==`Tzero & phi1)
			 | (OP==`JMP_abs & T==`Tone & phi1)
			 | (OP==`JMP_abs & T==`Ttwo & phi1)
			 | (OP==`EOR_abs & T==`Tzero & phi1)
			 | (OP==`EOR_abs & T==`Tone & phi1)
			 | (OP==`EOR_abs & T==`Ttwo & phi1)
			 | (OP==`EOR_abs & T==`Tthree & phi1)
			 | (OP==`LSR_abs & T==`Tzero & phi1)
			 | (OP==`LSR_abs & T==`Tone & phi1)
			 | (OP==`LSR_abs & T==`Ttwo & phi1)
			 | (OP==`LSR_abs & T==`Tthree & phi1)
			 | (OP==`LSR_abs & T==`Tfour & phi1)
			 | (OP==`LSR_abs & T==`Tfive & phi1)
			 | (OP==`BVC_rel & T==`Tzero & phi1)
			 | (OP==`BVC_rel & T==`Ttwo & phi1)
			 | (OP==`BVC_rel & T==`Tthree & phi1)
			 | (OP==`BVC_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BVC_rel & T==`T1BranchCross & phi1)
			 | (OP==`BVC_rel & T==`T1NoBranch & phi1)
			 | (OP==`EOR_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`EOR_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`EOR_izy & T==`Tone & phi1)
			 | (OP==`EOR_izy & T==`Ttwo & phi1)
			 | (OP==`EOR_izy & T==`Tthree & phi1)
			 | (OP==`EOR_izy & T==`Tfour & phi1)
			 | (OP==`EOR_izy & T==`Tfive & phi1)
			 | (OP==`EOR_zpx & T==`Tzero & phi1)
			 | (OP==`EOR_zpx & T==`Tone & phi1)
			 | (OP==`EOR_zpx & T==`Ttwo & phi1)
			 | (OP==`EOR_zpx & T==`Tthree & phi1)
			 | (OP==`LSR_zpx & T==`Tzero & phi1)
			 | (OP==`LSR_zpx & T==`Tone & phi1)
			 | (OP==`LSR_zpx & T==`Ttwo & phi1)
			 | (OP==`LSR_zpx & T==`Tthree & phi1)
			 | (OP==`LSR_zpx & T==`Tfour & phi1)
			 | (OP==`LSR_zpx & T==`Tfive & phi1)
			 | (OP==`CLI & T==`Tone & phi1)
			 | (OP==`CLI & T==`Ttwo & phi1)
			 | (OP==`EOR_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`EOR_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`EOR_aby & T==`Tone & phi1)
			 | (OP==`EOR_aby & T==`Ttwo & phi1)
			 | (OP==`EOR_aby & T==`Tthree & phi1)
			 | (OP==`EOR_aby & T==`Tfour & phi1)
			 | (OP==`EOR_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`EOR_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`EOR_abx & T==`Tone & phi1)
			 | (OP==`EOR_abx & T==`Ttwo & phi1)
			 | (OP==`EOR_abx & T==`Tthree & phi1)
			 | (OP==`EOR_abx & T==`Tfour & phi1)
			 | (OP==`LSR_abx & T==`Tzero & phi1)
			 | (OP==`LSR_abx & T==`Tone & phi1)
			 | (OP==`LSR_abx & T==`Ttwo & phi1)
			 | (OP==`LSR_abx & T==`Tthree & phi1)
			 | (OP==`LSR_abx & T==`Tfour & phi1)
			 | (OP==`LSR_abx & T==`Tfive & phi1)
			 | (OP==`LSR_abx & T==`Tsix & phi1)
			 | (OP==`RTS & T==`Tzero & phi1)
			 | (OP==`RTS & T==`Tone & phi1)
			 | (OP==`RTS & T==`Ttwo & phi1)
			 | (OP==`RTS & T==`Tthree & phi1)
			 | (OP==`RTS & T==`Tfour & phi1)
			 | (OP==`ADC_izx & T==`Tzero & phi1)
			 | (OP==`ADC_izx & T==`Tone & phi1)
			 | (OP==`ADC_izx & T==`Ttwo & phi1)
			 | (OP==`ADC_izx & T==`Tthree & phi1)
			 | (OP==`ADC_izx & T==`Tfour & phi1)
			 | (OP==`ADC_izx & T==`Tfive & phi1)
			 | (OP==`ADC_zp & T==`Tzero & phi1)
			 | (OP==`ADC_zp & T==`Tone & phi1)
			 | (OP==`ADC_zp & T==`Ttwo & phi1)
			 | (OP==`ROR_zp & T==`Tzero & phi1)
			 | (OP==`ROR_zp & T==`Tone & phi1)
			 | (OP==`ROR_zp & T==`Ttwo & phi1)
			 | (OP==`ROR_zp & T==`Tthree & phi1)
			 | (OP==`ROR_zp & T==`Tfour & phi1)
			 | (OP==`PLA & T==`Tone & phi1)
			 | (OP==`PLA & T==`Ttwo & phi1)
			 | (OP==`PLA & T==`Tthree & phi1)
			 | (OP==`ADC_imm & T==`Tone & phi1)
			 | (OP==`ADC_imm & T==`Ttwo & phi1)
			 | (OP==`ROR & T==`Tone & phi1)
			 | (OP==`ROR & T==`Ttwo & phi1)
			 | (OP==`JMP_zp & T==`Tzero & phi1)
			 | (OP==`JMP_zp & T==`Tone & phi1)
			 | (OP==`JMP_zp & T==`Ttwo & phi1)
			 | (OP==`JMP_zp & T==`Tthree & phi1)
			 | (OP==`JMP_zp & T==`Tfour & phi1)
			 | (OP==`ADC_abs & T==`Tzero & phi1)
			 | (OP==`ADC_abs & T==`Tone & phi1)
			 | (OP==`ADC_abs & T==`Ttwo & phi1)
			 | (OP==`ADC_abs & T==`Tthree & phi1)
			 | (OP==`ROR_abs & T==`Tzero & phi1)
			 | (OP==`ROR_abs & T==`Tone & phi1)
			 | (OP==`ROR_abs & T==`Ttwo & phi1)
			 | (OP==`ROR_abs & T==`Tthree & phi1)
			 | (OP==`ROR_abs & T==`Tfour & phi1)
			 | (OP==`ROR_abs & T==`Tfive & phi1)
			 | (OP==`BVS_rel & T==`Tzero & phi1)
			 | (OP==`BVS_rel & T==`Ttwo & phi1)
			 | (OP==`BVS_rel & T==`Tthree & phi1)
			 | (OP==`BVS_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BVS_rel & T==`T1BranchCross & phi1)
			 | (OP==`BVS_rel & T==`T1NoBranch & phi1)
			 | (OP==`ADC_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ADC_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`ADC_izy & T==`Tone & phi1)
			 | (OP==`ADC_izy & T==`Ttwo & phi1)
			 | (OP==`ADC_izy & T==`Tthree & phi1)
			 | (OP==`ADC_izy & T==`Tfour & phi1)
			 | (OP==`ADC_izy & T==`Tfive & phi1)
			 | (OP==`ADC_zpx & T==`Tzero & phi1)
			 | (OP==`ADC_zpx & T==`Tone & phi1)
			 | (OP==`ADC_zpx & T==`Ttwo & phi1)
			 | (OP==`ADC_zpx & T==`Tthree & phi1)
			 | (OP==`ROR_zpx & T==`Tzero & phi1)
			 | (OP==`ROR_zpx & T==`Tone & phi1)
			 | (OP==`ROR_zpx & T==`Ttwo & phi1)
			 | (OP==`ROR_zpx & T==`Tthree & phi1)
			 | (OP==`ROR_zpx & T==`Tfour & phi1)
			 | (OP==`ROR_zpx & T==`Tfive & phi1)
			 | (OP==`SEI & T==`Tone & phi1)
			 | (OP==`SEI & T==`Ttwo & phi1)
			 | (OP==`ADC_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ADC_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`ADC_aby & T==`Tone & phi1)
			 | (OP==`ADC_aby & T==`Ttwo & phi1)
			 | (OP==`ADC_aby & T==`Tthree & phi1)
			 | (OP==`ADC_aby & T==`Tfour & phi1)
			 | (OP==`ADC_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ADC_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`ADC_abx & T==`Tone & phi1)
			 | (OP==`ADC_abx & T==`Ttwo & phi1)
			 | (OP==`ADC_abx & T==`Tthree & phi1)
			 | (OP==`ADC_abx & T==`Tfour & phi1)
			 | (OP==`ROR_abx & T==`Tzero & phi1)
			 | (OP==`ROR_abx & T==`Tone & phi1)
			 | (OP==`ROR_abx & T==`Ttwo & phi1)
			 | (OP==`ROR_abx & T==`Tthree & phi1)
			 | (OP==`ROR_abx & T==`Tfour & phi1)
			 | (OP==`ROR_abx & T==`Tfive & phi1)
			 | (OP==`ROR_abx & T==`Tsix & phi1)
			 | (OP==`STA_izx & T==`Tzero & phi1)
			 | (OP==`STA_izx & T==`Tone & phi1)
			 | (OP==`STA_izx & T==`Ttwo & phi1)
			 | (OP==`STA_izx & T==`Tthree & phi1)
			 | (OP==`STA_izx & T==`Tfour & phi1)
			 | (OP==`STA_izx & T==`Tfive & phi1)
			 | (OP==`STY_zp & T==`Tzero & phi1)
			 | (OP==`STY_zp & T==`Tone & phi1)
			 | (OP==`STY_zp & T==`Ttwo & phi1)
			 | (OP==`STA_zp & T==`Tzero & phi1)
			 | (OP==`STA_zp & T==`Tone & phi1)
			 | (OP==`STA_zp & T==`Ttwo & phi1)
			 | (OP==`STX_zp & T==`Tzero & phi1)
			 | (OP==`STX_zp & T==`Tone & phi1)
			 | (OP==`STX_zp & T==`Ttwo & phi1)
			 | (OP==`DEY & T==`Tone & phi1)
			 | (OP==`DEY & T==`Ttwo & phi1)
			 | (OP==`TXA & T==`Tone & phi1)
			 | (OP==`TXA & T==`Ttwo & phi1)
			 | (OP==`STY_abs & T==`Tzero & phi1)
			 | (OP==`STY_abs & T==`Tone & phi1)
			 | (OP==`STY_abs & T==`Ttwo & phi1)
			 | (OP==`STY_abs & T==`Tthree & phi1)
			 | (OP==`STA_abs & T==`Tzero & phi1)
			 | (OP==`STA_abs & T==`Tone & phi1)
			 | (OP==`STA_abs & T==`Ttwo & phi1)
			 | (OP==`STA_abs & T==`Tthree & phi1)
			 | (OP==`STX_abs & T==`Tzero & phi1)
			 | (OP==`STX_abs & T==`Tone & phi1)
			 | (OP==`STX_abs & T==`Ttwo & phi1)
			 | (OP==`STX_abs & T==`Tthree & phi1)
			 | (OP==`BCC_rel & T==`Tzero & phi1)
			 | (OP==`BCC_rel & T==`Ttwo & phi1)
			 | (OP==`BCC_rel & T==`Tthree & phi1)
			 | (OP==`BCC_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BCC_rel & T==`T1BranchCross & phi1)
			 | (OP==`BCC_rel & T==`T1NoBranch & phi1)
			 | (OP==`STA_izy & T==`Tzero & phi1)
			 | (OP==`STA_izy & T==`Tone & phi1)
			 | (OP==`STA_izy & T==`Ttwo & phi1)
			 | (OP==`STA_izy & T==`Tthree & phi1)
			 | (OP==`STA_izy & T==`Tfour & phi1)
			 | (OP==`STA_izy & T==`Tfive & phi1)
			 | (OP==`STY_zpx & T==`Tzero & phi1)
			 | (OP==`STY_zpx & T==`Tone & phi1)
			 | (OP==`STY_zpx & T==`Ttwo & phi1)
			 | (OP==`STY_zpx & T==`Tthree & phi1)
			 | (OP==`STA_zpx & T==`Tzero & phi1)
			 | (OP==`STA_zpx & T==`Tone & phi1)
			 | (OP==`STA_zpx & T==`Ttwo & phi1)
			 | (OP==`STA_zpx & T==`Tthree & phi1)
			 | (OP==`STX_zpy & T==`Tzero & phi1)
			 | (OP==`STX_zpy & T==`Tone & phi1)
			 | (OP==`STX_zpy & T==`Ttwo & phi1)
			 | (OP==`STX_zpy & T==`Tthree & phi1)
			 | (OP==`TYA & T==`Tone & phi1)
			 | (OP==`TYA & T==`Ttwo & phi1)
			 | (OP==`STA_aby & T==`Tzero & phi1)
			 | (OP==`STA_aby & T==`Tone & phi1)
			 | (OP==`STA_aby & T==`Ttwo & phi1)
			 | (OP==`STA_aby & T==`Tthree & phi1)
			 | (OP==`STA_aby & T==`Tfour & phi1)
			 | (OP==`TXS & T==`Ttwo & phi1)
			 | (OP==`STA_abx & T==`Tzero & phi1)
			 | (OP==`STA_abx & T==`Tone & phi1)
			 | (OP==`STA_abx & T==`Ttwo & phi1)
			 | (OP==`STA_abx & T==`Tthree & phi1)
			 | (OP==`STA_abx & T==`Tfour & phi1)
			 | (OP==`LDY_imm & T==`Tone & phi1)
			 | (OP==`LDY_imm & T==`Ttwo & phi1)
			 | (OP==`LDA_izx & T==`Tzero & phi1)
			 | (OP==`LDA_izx & T==`Tone & phi1)
			 | (OP==`LDA_izx & T==`Ttwo & phi1)
			 | (OP==`LDA_izx & T==`Tthree & phi1)
			 | (OP==`LDA_izx & T==`Tfour & phi1)
			 | (OP==`LDA_izx & T==`Tfive & phi1)
			 | (OP==`LDX_imm & T==`Tone & phi1)
			 | (OP==`LDX_imm & T==`Ttwo & phi1)
			 | (OP==`LDY_zp & T==`Tzero & phi1)
			 | (OP==`LDY_zp & T==`Tone & phi1)
			 | (OP==`LDY_zp & T==`Ttwo & phi1)
			 | (OP==`LDA_zp & T==`Tzero & phi1)
			 | (OP==`LDA_zp & T==`Tone & phi1)
			 | (OP==`LDA_zp & T==`Ttwo & phi1)
			 | (OP==`LDX_zp & T==`Tzero & phi1)
			 | (OP==`LDX_zp & T==`Tone & phi1)
			 | (OP==`LDX_zp & T==`Ttwo & phi1)
			 | (OP==`TAY & T==`Tone & phi1)
			 | (OP==`TAY & T==`Ttwo & phi1)
			 | (OP==`LDA_imm & T==`Tone & phi1)
			 | (OP==`LDA_imm & T==`Ttwo & phi1)
			 | (OP==`TAX & T==`Tone & phi1)
			 | (OP==`TAX & T==`Ttwo & phi1)
			 | (OP==`LDY_abs & T==`Tzero & phi1)
			 | (OP==`LDY_abs & T==`Tone & phi1)
			 | (OP==`LDY_abs & T==`Ttwo & phi1)
			 | (OP==`LDY_abs & T==`Tthree & phi1)
			 | (OP==`LDA_abs & T==`Tzero & phi1)
			 | (OP==`LDA_abs & T==`Tone & phi1)
			 | (OP==`LDA_abs & T==`Ttwo & phi1)
			 | (OP==`LDA_abs & T==`Tthree & phi1)
			 | (OP==`LDX_abs & T==`Tzero & phi1)
			 | (OP==`LDX_abs & T==`Tone & phi1)
			 | (OP==`LDX_abs & T==`Ttwo & phi1)
			 | (OP==`LDX_abs & T==`Tthree & phi1)
			 | (OP==`BCS_rel & T==`Tzero & phi1)
			 | (OP==`BCS_rel & T==`Ttwo & phi1)
			 | (OP==`BCS_rel & T==`Tthree & phi1)
			 | (OP==`BCS_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BCS_rel & T==`T1BranchCross & phi1)
			 | (OP==`BCS_rel & T==`T1NoBranch & phi1)
			 | (OP==`LDA_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDA_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`LDA_izy & T==`Tone & phi1)
			 | (OP==`LDA_izy & T==`Ttwo & phi1)
			 | (OP==`LDA_izy & T==`Tthree & phi1)
			 | (OP==`LDA_izy & T==`Tfour & phi1)
			 | (OP==`LDA_izy & T==`Tfive & phi1)
			 | (OP==`LDY_zpx & T==`Tzero & phi1)
			 | (OP==`LDY_zpx & T==`Tone & phi1)
			 | (OP==`LDY_zpx & T==`Ttwo & phi1)
			 | (OP==`LDY_zpx & T==`Tthree & phi1)
			 | (OP==`LDA_zpx & T==`Tzero & phi1)
			 | (OP==`LDA_zpx & T==`Tone & phi1)
			 | (OP==`LDA_zpx & T==`Ttwo & phi1)
			 | (OP==`LDA_zpx & T==`Tthree & phi1)
			 | (OP==`LDX_zpy & T==`Tzero & phi1)
			 | (OP==`LDX_zpy & T==`Tone & phi1)
			 | (OP==`LDX_zpy & T==`Ttwo & phi1)
			 | (OP==`LDX_zpy & T==`Tthree & phi1)
			 | (OP==`CLV & T==`Tone & phi1)
			 | (OP==`CLV & T==`Ttwo & phi1)
			 | (OP==`LDA_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDA_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`LDA_aby & T==`Tone & phi1)
			 | (OP==`LDA_aby & T==`Ttwo & phi1)
			 | (OP==`LDA_aby & T==`Tthree & phi1)
			 | (OP==`LDA_aby & T==`Tfour & phi1)
			 | (OP==`TSX & T==`Tone & phi1)
			 | (OP==`TSX & T==`Ttwo & phi1)
			 | (OP==`LDY_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDY_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`LDY_abx & T==`Tone & phi1)
			 | (OP==`LDY_abx & T==`Ttwo & phi1)
			 | (OP==`LDY_abx & T==`Tthree & phi1)
			 | (OP==`LDY_abx & T==`Tfour & phi1)
			 | (OP==`LDA_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDA_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`LDA_abx & T==`Tone & phi1)
			 | (OP==`LDA_abx & T==`Ttwo & phi1)
			 | (OP==`LDA_abx & T==`Tthree & phi1)
			 | (OP==`LDA_abx & T==`Tfour & phi1)
			 | (OP==`LDX_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDX_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`LDX_aby & T==`Tone & phi1)
			 | (OP==`LDX_aby & T==`Ttwo & phi1)
			 | (OP==`LDX_aby & T==`Tthree & phi1)
			 | (OP==`LDX_aby & T==`Tfour & phi1)
			 | (OP==`CPY_imm & T==`Tone & phi1)
			 | (OP==`CPY_imm & T==`Ttwo & phi1)
			 | (OP==`CMP_izx & T==`Tzero & phi1)
			 | (OP==`CMP_izx & T==`Tone & phi1)
			 | (OP==`CMP_izx & T==`Ttwo & phi1)
			 | (OP==`CMP_izx & T==`Tthree & phi1)
			 | (OP==`CMP_izx & T==`Tfour & phi1)
			 | (OP==`CMP_izx & T==`Tfive & phi1)
			 | (OP==`CPY_zp & T==`Tzero & phi1)
			 | (OP==`CPY_zp & T==`Tone & phi1)
			 | (OP==`CPY_zp & T==`Ttwo & phi1)
			 | (OP==`CMP_zp & T==`Tzero & phi1)
			 | (OP==`CMP_zp & T==`Tone & phi1)
			 | (OP==`CMP_zp & T==`Ttwo & phi1)
			 | (OP==`DEC_zp & T==`Tzero & phi1)
			 | (OP==`DEC_zp & T==`Tone & phi1)
			 | (OP==`DEC_zp & T==`Ttwo & phi1)
			 | (OP==`DEC_zp & T==`Tthree & phi1)
			 | (OP==`DEC_zp & T==`Tfour & phi1)
			 | (OP==`INY & T==`Tone & phi1)
			 | (OP==`INY & T==`Ttwo & phi1)
			 | (OP==`CMP_imm & T==`Tone & phi1)
			 | (OP==`CMP_imm & T==`Ttwo & phi1)
			 | (OP==`DEX & T==`Tone & phi1)
			 | (OP==`DEX & T==`Ttwo & phi1)
			 | (OP==`CPY_abs & T==`Tzero & phi1)
			 | (OP==`CPY_abs & T==`Tone & phi1)
			 | (OP==`CPY_abs & T==`Ttwo & phi1)
			 | (OP==`CPY_abs & T==`Tthree & phi1)
			 | (OP==`CMP_abs & T==`Tzero & phi1)
			 | (OP==`CMP_abs & T==`Tone & phi1)
			 | (OP==`CMP_abs & T==`Ttwo & phi1)
			 | (OP==`CMP_abs & T==`Tthree & phi1)
			 | (OP==`DEC_abs & T==`Tzero & phi1)
			 | (OP==`DEC_abs & T==`Tone & phi1)
			 | (OP==`DEC_abs & T==`Ttwo & phi1)
			 | (OP==`DEC_abs & T==`Tthree & phi1)
			 | (OP==`DEC_abs & T==`Tfour & phi1)
			 | (OP==`DEC_abs & T==`Tfive & phi1)
			 | (OP==`BNE_rel & T==`Tzero & phi1)
			 | (OP==`BNE_rel & T==`Ttwo & phi1)
			 | (OP==`BNE_rel & T==`Tthree & phi1)
			 | (OP==`BNE_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BNE_rel & T==`T1BranchCross & phi1)
			 | (OP==`BNE_rel & T==`T1NoBranch & phi1)
			 | (OP==`CMP_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`CMP_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`CMP_izy & T==`Tone & phi1)
			 | (OP==`CMP_izy & T==`Ttwo & phi1)
			 | (OP==`CMP_izy & T==`Tthree & phi1)
			 | (OP==`CMP_izy & T==`Tfour & phi1)
			 | (OP==`CMP_izy & T==`Tfive & phi1)
			 | (OP==`CMP_zpx & T==`Tzero & phi1)
			 | (OP==`CMP_zpx & T==`Tone & phi1)
			 | (OP==`CMP_zpx & T==`Ttwo & phi1)
			 | (OP==`CMP_zpx & T==`Tthree & phi1)
			 | (OP==`DEC_zpx & T==`Tzero & phi1)
			 | (OP==`DEC_zpx & T==`Tone & phi1)
			 | (OP==`DEC_zpx & T==`Ttwo & phi1)
			 | (OP==`DEC_zpx & T==`Tthree & phi1)
			 | (OP==`DEC_zpx & T==`Tfour & phi1)
			 | (OP==`DEC_zpx & T==`Tfive & phi1)
			 | (OP==`CLD & T==`Tone & phi1)
			 | (OP==`CLD & T==`Ttwo & phi1)
			 | (OP==`CMP_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`CMP_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`CMP_aby & T==`Tone & phi1)
			 | (OP==`CMP_aby & T==`Ttwo & phi1)
			 | (OP==`CMP_aby & T==`Tthree & phi1)
			 | (OP==`CMP_aby & T==`Tfour & phi1)
			 | (OP==`CMP_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`CMP_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`CMP_abx & T==`Tone & phi1)
			 | (OP==`CMP_abx & T==`Ttwo & phi1)
			 | (OP==`CMP_abx & T==`Tthree & phi1)
			 | (OP==`CMP_abx & T==`Tfour & phi1)
			 | (OP==`DEC_abx & T==`Tzero & phi1)
			 | (OP==`DEC_abx & T==`Tone & phi1)
			 | (OP==`DEC_abx & T==`Ttwo & phi1)
			 | (OP==`DEC_abx & T==`Tthree & phi1)
			 | (OP==`DEC_abx & T==`Tfour & phi1)
			 | (OP==`DEC_abx & T==`Tfive & phi1)
			 | (OP==`DEC_abx & T==`Tsix & phi1)
			 | (OP==`CPX_imm & T==`Tone & phi1)
			 | (OP==`CPX_imm & T==`Ttwo & phi1)
			 | (OP==`SBC_izx & T==`Tzero & phi1)
			 | (OP==`SBC_izx & T==`Tone & phi1)
			 | (OP==`SBC_izx & T==`Ttwo & phi1)
			 | (OP==`SBC_izx & T==`Tthree & phi1)
			 | (OP==`SBC_izx & T==`Tfour & phi1)
			 | (OP==`SBC_izx & T==`Tfive & phi1)
			 | (OP==`CPX_zp & T==`Tzero & phi1)
			 | (OP==`CPX_zp & T==`Tone & phi1)
			 | (OP==`CPX_zp & T==`Ttwo & phi1)
			 | (OP==`SBC_zp & T==`Tzero & phi1)
			 | (OP==`SBC_zp & T==`Tone & phi1)
			 | (OP==`SBC_zp & T==`Ttwo & phi1)
			 | (OP==`INC_zp & T==`Tzero & phi1)
			 | (OP==`INC_zp & T==`Tone & phi1)
			 | (OP==`INC_zp & T==`Ttwo & phi1)
			 | (OP==`INC_zp & T==`Tthree & phi1)
			 | (OP==`INC_zp & T==`Tfour & phi1)
			 | (OP==`INX & T==`Tone & phi1)
			 | (OP==`INX & T==`Ttwo & phi1)
			 | (OP==`SBC_imm & T==`Tone & phi1)
			 | (OP==`SBC_imm & T==`Ttwo & phi1)
			 | (OP==`NOP & T==`Tone & phi1)
			 | (OP==`NOP & T==`Ttwo & phi1)
			 | (OP==`CPX_abs & T==`Tzero & phi1)
			 | (OP==`CPX_abs & T==`Tone & phi1)
			 | (OP==`CPX_abs & T==`Ttwo & phi1)
			 | (OP==`CPX_abs & T==`Tthree & phi1)
			 | (OP==`SBC_abs & T==`Tzero & phi1)
			 | (OP==`SBC_abs & T==`Tone & phi1)
			 | (OP==`SBC_abs & T==`Ttwo & phi1)
			 | (OP==`SBC_abs & T==`Tthree & phi1)
			 | (OP==`INC_abs & T==`Tzero & phi1)
			 | (OP==`INC_abs & T==`Tone & phi1)
			 | (OP==`INC_abs & T==`Ttwo & phi1)
			 | (OP==`INC_abs & T==`Tthree & phi1)
			 | (OP==`INC_abs & T==`Tfour & phi1)
			 | (OP==`INC_abs & T==`Tfive & phi1)
			 | (OP==`BEQ_rel & T==`Tzero & phi1)
			 | (OP==`BEQ_rel & T==`Ttwo & phi1)
			 | (OP==`BEQ_rel & T==`Tthree & phi1)
			 | (OP==`BEQ_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BEQ_rel & T==`T1BranchCross & phi1)
			 | (OP==`BEQ_rel & T==`T1NoBranch & phi1)
			 | (OP==`SBC_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`SBC_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`SBC_izy & T==`Tone & phi1)
			 | (OP==`SBC_izy & T==`Ttwo & phi1)
			 | (OP==`SBC_izy & T==`Tthree & phi1)
			 | (OP==`SBC_izy & T==`Tfour & phi1)
			 | (OP==`SBC_izy & T==`Tfive & phi1)
			 | (OP==`SBC_zpx & T==`Tzero & phi1)
			 | (OP==`SBC_zpx & T==`Tone & phi1)
			 | (OP==`SBC_zpx & T==`Ttwo & phi1)
			 | (OP==`SBC_zpx & T==`Tthree & phi1)
			 | (OP==`INC_zpx & T==`Tzero & phi1)
			 | (OP==`INC_zpx & T==`Tone & phi1)
			 | (OP==`INC_zpx & T==`Ttwo & phi1)
			 | (OP==`INC_zpx & T==`Tthree & phi1)
			 | (OP==`INC_zpx & T==`Tfour & phi1)
			 | (OP==`INC_zpx & T==`Tfive & phi1)
			 | (OP==`SED & T==`Tone & phi1)
			 | (OP==`SED & T==`Ttwo & phi1)
			 | (OP==`SBC_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`SBC_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`SBC_aby & T==`Tone & phi1)
			 | (OP==`SBC_aby & T==`Ttwo & phi1)
			 | (OP==`SBC_aby & T==`Tthree & phi1)
			 | (OP==`SBC_aby & T==`Tfour & phi1)
			 | (OP==`SBC_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`SBC_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`SBC_abx & T==`Tone & phi1)
			 | (OP==`SBC_abx & T==`Ttwo & phi1)
			 | (OP==`SBC_abx & T==`Tthree & phi1)
			 | (OP==`SBC_abx & T==`Tfour & phi1)
			 | (OP==`INC_abx & T==`Tzero & phi1)
			 | (OP==`INC_abx & T==`Tone & phi1)
			 | (OP==`INC_abx & T==`Ttwo & phi1)
			 | (OP==`INC_abx & T==`Tthree & phi1)
			 | (OP==`INC_abx & T==`Tfour & phi1)
			 | (OP==`INC_abx & T==`Tfive & phi1)
			 | (OP==`INC_abx & T==`Tsix & phi1)
			;

assign control[`S_SB] = (OP==`TSX & T==`Tone & phi1)
			 | (OP==`TSX & T==`Ttwo & phi2)
			;

assign control[`DB_L_ADD] = (OP==`BPL_rel & T==`Tzero & phi1)
			 | (OP==`BPL_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`JSR_abs & T==`Tzero & phi1)
			 | (OP==`BMI_rel & T==`Tzero & phi1)
			 | (OP==`BMI_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BVC_rel & T==`Tzero & phi1)
			 | (OP==`BVC_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BVS_rel & T==`Tzero & phi1)
			 | (OP==`BVS_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BCC_rel & T==`Tzero & phi1)
			 | (OP==`BCC_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BCS_rel & T==`Tzero & phi1)
			 | (OP==`BCS_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`CPY_imm & T==`Tone & phi1)
			 | (OP==`CMP_izx & T==`Tone & phi1)
			 | (OP==`CPY_zp & T==`Tone & phi1)
			 | (OP==`CMP_zp & T==`Tone & phi1)
			 | (OP==`INY & T==`Tone & phi1)
			 | (OP==`CMP_imm & T==`Tone & phi1)
			 | (OP==`CPY_abs & T==`Tone & phi1)
			 | (OP==`CMP_abs & T==`Tone & phi1)
			 | (OP==`BNE_rel & T==`Tzero & phi1)
			 | (OP==`BNE_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`CMP_izy & T==`Tone & phi1)
			 | (OP==`CMP_zpx & T==`Tone & phi1)
			 | (OP==`CMP_aby & T==`Tone & phi1)
			 | (OP==`CMP_abx & T==`Tone & phi1)
			 | (OP==`CPX_imm & T==`Tone & phi1)
			 | (OP==`SBC_izx & T==`Tone & phi1)
			 | (OP==`CPX_zp & T==`Tone & phi1)
			 | (OP==`SBC_zp & T==`Tone & phi1)
			 | (OP==`INX & T==`Tone & phi1)
			 | (OP==`SBC_imm & T==`Tone & phi1)
			 | (OP==`CPX_abs & T==`Tone & phi1)
			 | (OP==`SBC_abs & T==`Tone & phi1)
			 | (OP==`BEQ_rel & T==`Tzero & phi1)
			 | (OP==`BEQ_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`SBC_izy & T==`Tone & phi1)
			 | (OP==`SBC_zpx & T==`Tone & phi1)
			 | (OP==`SBC_aby & T==`Tone & phi1)
			 | (OP==`SBC_abx & T==`Tone & phi1)
			;

assign control[`DB_ADD] = (OP==`BRK & T==`Tzero & phi1)
			 | (OP==`BRK & T==`Tone & phi1)
			 | (OP==`BRK & T==`Ttwo & phi1)
			 | (OP==`BRK & T==`Tsix & phi1)
			 | (OP==`ORA_izx & T==`Tzero & phi1)
			 | (OP==`ORA_izx & T==`Tone & phi1)
			 | (OP==`ORA_izx & T==`Ttwo & phi1)
			 | (OP==`ORA_izx & T==`Tfive & phi1)
			 | (OP==`ORA_zp & T==`Tone & phi1)
			 | (OP==`ORA_zp & T==`Ttwo & phi1)
			 | (OP==`ASL_zp & T==`Tzero & phi1)
			 | (OP==`ASL_zp & T==`Tone & phi1)
			 | (OP==`ASL_zp & T==`Ttwo & phi1)
			 | (OP==`ASL_zp & T==`Tfour & phi1)
			 | (OP==`PHP & T==`Tone & phi1)
			 | (OP==`PHP & T==`Ttwo & phi1)
			 | (OP==`ORA_imm & T==`Tone & phi1)
			 | (OP==`ORA_imm & T==`Ttwo & phi1)
			 | (OP==`ASL & T==`Tone & phi1)
			 | (OP==`ASL & T==`Ttwo & phi1)
			 | (OP==`ORA_abs & T==`Tzero & phi1)
			 | (OP==`ORA_abs & T==`Tone & phi1)
			 | (OP==`ORA_abs & T==`Ttwo & phi1)
			 | (OP==`ORA_abs & T==`Tthree & phi1)
			 | (OP==`ASL_abs & T==`Tzero & phi1)
			 | (OP==`ASL_abs & T==`Tone & phi1)
			 | (OP==`ASL_abs & T==`Ttwo & phi1)
			 | (OP==`ASL_abs & T==`Tthree & phi1)
			 | (OP==`ASL_abs & T==`Tfour & phi1)
			 | (OP==`ASL_abs & T==`Tfive & phi1)
			 | (OP==`BPL_rel & T==`Ttwo & phi1)
			 | (OP==`BPL_rel & T==`T1BranchCross & phi1)
			 | (OP==`ORA_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`ORA_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ORA_izy & T==`Tone & phi1)
			 | (OP==`ORA_izy & T==`Ttwo & phi1)
			 | (OP==`ORA_izy & T==`Tfour & phi1)
			 | (OP==`ORA_izy & T==`Tfive & phi1)
			 | (OP==`ORA_zpx & T==`Tzero & phi1)
			 | (OP==`ORA_zpx & T==`Tone & phi1)
			 | (OP==`ORA_zpx & T==`Ttwo & phi1)
			 | (OP==`ASL_zpx & T==`Tzero & phi1)
			 | (OP==`ASL_zpx & T==`Tone & phi1)
			 | (OP==`ASL_zpx & T==`Ttwo & phi1)
			 | (OP==`ASL_zpx & T==`Tfour & phi1)
			 | (OP==`ASL_zpx & T==`Tfive & phi1)
			 | (OP==`CLC & T==`Tone & phi1)
			 | (OP==`CLC & T==`Ttwo & phi1)
			 | (OP==`ORA_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ORA_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`ORA_aby & T==`Tone & phi1)
			 | (OP==`ORA_aby & T==`Ttwo & phi1)
			 | (OP==`ORA_aby & T==`Tthree & phi1)
			 | (OP==`ORA_aby & T==`Tfour & phi1)
			 | (OP==`ORA_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ORA_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`ORA_abx & T==`Tone & phi1)
			 | (OP==`ORA_abx & T==`Ttwo & phi1)
			 | (OP==`ORA_abx & T==`Tthree & phi1)
			 | (OP==`ORA_abx & T==`Tfour & phi1)
			 | (OP==`ASL_abx & T==`Tzero & phi1)
			 | (OP==`ASL_abx & T==`Tone & phi1)
			 | (OP==`ASL_abx & T==`Ttwo & phi1)
			 | (OP==`ASL_abx & T==`Tthree & phi1)
			 | (OP==`ASL_abx & T==`Tfour & phi1)
			 | (OP==`ASL_abx & T==`Tfive & phi1)
			 | (OP==`ASL_abx & T==`Tsix & phi1)
			 | (OP==`JSR_abs & T==`Tone & phi1)
			 | (OP==`JSR_abs & T==`Ttwo & phi1)
			 | (OP==`AND_izx & T==`Tzero & phi1)
			 | (OP==`AND_izx & T==`Tone & phi1)
			 | (OP==`AND_izx & T==`Ttwo & phi1)
			 | (OP==`AND_izx & T==`Tfive & phi1)
			 | (OP==`BIT_zp & T==`Tone & phi1)
			 | (OP==`BIT_zp & T==`Ttwo & phi1)
			 | (OP==`AND_zp & T==`Tone & phi1)
			 | (OP==`AND_zp & T==`Ttwo & phi1)
			 | (OP==`ROL_zp & T==`Tzero & phi1)
			 | (OP==`ROL_zp & T==`Tone & phi1)
			 | (OP==`ROL_zp & T==`Ttwo & phi1)
			 | (OP==`ROL_zp & T==`Tfour & phi1)
			 | (OP==`PLP & T==`Tone & phi1)
			 | (OP==`PLP & T==`Ttwo & phi1)
			 | (OP==`AND_imm & T==`Tone & phi1)
			 | (OP==`AND_imm & T==`Ttwo & phi1)
			 | (OP==`ROL & T==`Tone & phi1)
			 | (OP==`ROL & T==`Ttwo & phi1)
			 | (OP==`BIT_abs & T==`Tone & phi1)
			 | (OP==`BIT_abs & T==`Ttwo & phi1)
			 | (OP==`BIT_abs & T==`Tthree & phi1)
			 | (OP==`AND_abs & T==`Tzero & phi1)
			 | (OP==`AND_abs & T==`Tone & phi1)
			 | (OP==`AND_abs & T==`Ttwo & phi1)
			 | (OP==`AND_abs & T==`Tthree & phi1)
			 | (OP==`ROL_abs & T==`Tzero & phi1)
			 | (OP==`ROL_abs & T==`Tone & phi1)
			 | (OP==`ROL_abs & T==`Ttwo & phi1)
			 | (OP==`ROL_abs & T==`Tthree & phi1)
			 | (OP==`ROL_abs & T==`Tfour & phi1)
			 | (OP==`ROL_abs & T==`Tfive & phi1)
			 | (OP==`BMI_rel & T==`Ttwo & phi1)
			 | (OP==`BMI_rel & T==`T1BranchCross & phi1)
			 | (OP==`AND_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`AND_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`AND_izy & T==`Tone & phi1)
			 | (OP==`AND_izy & T==`Ttwo & phi1)
			 | (OP==`AND_izy & T==`Tfour & phi1)
			 | (OP==`AND_izy & T==`Tfive & phi1)
			 | (OP==`AND_zpx & T==`Tzero & phi1)
			 | (OP==`AND_zpx & T==`Tone & phi1)
			 | (OP==`AND_zpx & T==`Ttwo & phi1)
			 | (OP==`ROL_zpx & T==`Tzero & phi1)
			 | (OP==`ROL_zpx & T==`Tone & phi1)
			 | (OP==`ROL_zpx & T==`Ttwo & phi1)
			 | (OP==`ROL_zpx & T==`Tfour & phi1)
			 | (OP==`ROL_zpx & T==`Tfive & phi1)
			 | (OP==`SEC & T==`Tone & phi1)
			 | (OP==`SEC & T==`Ttwo & phi1)
			 | (OP==`AND_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`AND_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`AND_aby & T==`Tone & phi1)
			 | (OP==`AND_aby & T==`Ttwo & phi1)
			 | (OP==`AND_aby & T==`Tthree & phi1)
			 | (OP==`AND_aby & T==`Tfour & phi1)
			 | (OP==`AND_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`AND_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`AND_abx & T==`Tone & phi1)
			 | (OP==`AND_abx & T==`Ttwo & phi1)
			 | (OP==`AND_abx & T==`Tthree & phi1)
			 | (OP==`AND_abx & T==`Tfour & phi1)
			 | (OP==`ROL_abx & T==`Tzero & phi1)
			 | (OP==`ROL_abx & T==`Tone & phi1)
			 | (OP==`ROL_abx & T==`Ttwo & phi1)
			 | (OP==`ROL_abx & T==`Tthree & phi1)
			 | (OP==`ROL_abx & T==`Tfour & phi1)
			 | (OP==`ROL_abx & T==`Tfive & phi1)
			 | (OP==`ROL_abx & T==`Tsix & phi1)
			 | (OP==`RTI & T==`Tzero & phi1)
			 | (OP==`RTI & T==`Tone & phi1)
			 | (OP==`RTI & T==`Ttwo & phi1)
			 | (OP==`EOR_izx & T==`Tzero & phi1)
			 | (OP==`EOR_izx & T==`Tone & phi1)
			 | (OP==`EOR_izx & T==`Ttwo & phi1)
			 | (OP==`EOR_izx & T==`Tfive & phi1)
			 | (OP==`EOR_zp & T==`Tone & phi1)
			 | (OP==`EOR_zp & T==`Ttwo & phi1)
			 | (OP==`LSR_zp & T==`Tzero & phi1)
			 | (OP==`LSR_zp & T==`Tone & phi1)
			 | (OP==`LSR_zp & T==`Ttwo & phi1)
			 | (OP==`LSR_zp & T==`Tfour & phi1)
			 | (OP==`PHA & T==`Tone & phi1)
			 | (OP==`PHA & T==`Ttwo & phi1)
			 | (OP==`EOR_imm & T==`Tone & phi1)
			 | (OP==`EOR_imm & T==`Ttwo & phi1)
			 | (OP==`LSR & T==`Tone & phi1)
			 | (OP==`LSR & T==`Ttwo & phi1)
			 | (OP==`JMP_abs & T==`Tzero & phi1)
			 | (OP==`JMP_abs & T==`Tone & phi1)
			 | (OP==`JMP_abs & T==`Ttwo & phi1)
			 | (OP==`EOR_abs & T==`Tzero & phi1)
			 | (OP==`EOR_abs & T==`Tone & phi1)
			 | (OP==`EOR_abs & T==`Ttwo & phi1)
			 | (OP==`EOR_abs & T==`Tthree & phi1)
			 | (OP==`LSR_abs & T==`Tzero & phi1)
			 | (OP==`LSR_abs & T==`Tone & phi1)
			 | (OP==`LSR_abs & T==`Ttwo & phi1)
			 | (OP==`LSR_abs & T==`Tthree & phi1)
			 | (OP==`LSR_abs & T==`Tfour & phi1)
			 | (OP==`LSR_abs & T==`Tfive & phi1)
			 | (OP==`BVC_rel & T==`Ttwo & phi1)
			 | (OP==`BVC_rel & T==`T1BranchCross & phi1)
			 | (OP==`EOR_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`EOR_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`EOR_izy & T==`Tone & phi1)
			 | (OP==`EOR_izy & T==`Ttwo & phi1)
			 | (OP==`EOR_izy & T==`Tfour & phi1)
			 | (OP==`EOR_izy & T==`Tfive & phi1)
			 | (OP==`EOR_zpx & T==`Tzero & phi1)
			 | (OP==`EOR_zpx & T==`Tone & phi1)
			 | (OP==`EOR_zpx & T==`Ttwo & phi1)
			 | (OP==`LSR_zpx & T==`Tzero & phi1)
			 | (OP==`LSR_zpx & T==`Tone & phi1)
			 | (OP==`LSR_zpx & T==`Ttwo & phi1)
			 | (OP==`LSR_zpx & T==`Tfour & phi1)
			 | (OP==`LSR_zpx & T==`Tfive & phi1)
			 | (OP==`CLI & T==`Tone & phi1)
			 | (OP==`CLI & T==`Ttwo & phi1)
			 | (OP==`EOR_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`EOR_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`EOR_aby & T==`Tone & phi1)
			 | (OP==`EOR_aby & T==`Ttwo & phi1)
			 | (OP==`EOR_aby & T==`Tthree & phi1)
			 | (OP==`EOR_aby & T==`Tfour & phi1)
			 | (OP==`EOR_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`EOR_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`EOR_abx & T==`Tone & phi1)
			 | (OP==`EOR_abx & T==`Ttwo & phi1)
			 | (OP==`EOR_abx & T==`Tthree & phi1)
			 | (OP==`EOR_abx & T==`Tfour & phi1)
			 | (OP==`LSR_abx & T==`Tzero & phi1)
			 | (OP==`LSR_abx & T==`Tone & phi1)
			 | (OP==`LSR_abx & T==`Ttwo & phi1)
			 | (OP==`LSR_abx & T==`Tthree & phi1)
			 | (OP==`LSR_abx & T==`Tfour & phi1)
			 | (OP==`LSR_abx & T==`Tfive & phi1)
			 | (OP==`LSR_abx & T==`Tsix & phi1)
			 | (OP==`RTS & T==`Tzero & phi1)
			 | (OP==`RTS & T==`Tone & phi1)
			 | (OP==`RTS & T==`Ttwo & phi1)
			 | (OP==`RTS & T==`Tfive & phi1)
			 | (OP==`ADC_izx & T==`Tzero & phi1)
			 | (OP==`ADC_izx & T==`Tone & phi1)
			 | (OP==`ADC_izx & T==`Ttwo & phi1)
			 | (OP==`ADC_izx & T==`Tfive & phi1)
			 | (OP==`ADC_zp & T==`Tone & phi1)
			 | (OP==`ADC_zp & T==`Ttwo & phi1)
			 | (OP==`ROR_zp & T==`Tzero & phi1)
			 | (OP==`ROR_zp & T==`Tone & phi1)
			 | (OP==`ROR_zp & T==`Ttwo & phi1)
			 | (OP==`ROR_zp & T==`Tfour & phi1)
			 | (OP==`PLA & T==`Tone & phi1)
			 | (OP==`PLA & T==`Ttwo & phi1)
			 | (OP==`ADC_imm & T==`Tone & phi1)
			 | (OP==`ADC_imm & T==`Ttwo & phi1)
			 | (OP==`ROR & T==`Tone & phi1)
			 | (OP==`ROR & T==`Ttwo & phi1)
			 | (OP==`JMP_zp & T==`Tzero & phi1)
			 | (OP==`JMP_zp & T==`Tone & phi1)
			 | (OP==`JMP_zp & T==`Ttwo & phi1)
			 | (OP==`JMP_zp & T==`Tthree & phi1)
			 | (OP==`ADC_abs & T==`Tzero & phi1)
			 | (OP==`ADC_abs & T==`Tone & phi1)
			 | (OP==`ADC_abs & T==`Ttwo & phi1)
			 | (OP==`ADC_abs & T==`Tthree & phi1)
			 | (OP==`ROR_abs & T==`Tzero & phi1)
			 | (OP==`ROR_abs & T==`Tone & phi1)
			 | (OP==`ROR_abs & T==`Ttwo & phi1)
			 | (OP==`ROR_abs & T==`Tthree & phi1)
			 | (OP==`ROR_abs & T==`Tfour & phi1)
			 | (OP==`ROR_abs & T==`Tfive & phi1)
			 | (OP==`BVS_rel & T==`Ttwo & phi1)
			 | (OP==`BVS_rel & T==`T1BranchCross & phi1)
			 | (OP==`ADC_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ADC_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`ADC_izy & T==`Tone & phi1)
			 | (OP==`ADC_izy & T==`Ttwo & phi1)
			 | (OP==`ADC_izy & T==`Tfour & phi1)
			 | (OP==`ADC_izy & T==`Tfive & phi1)
			 | (OP==`ADC_zpx & T==`Tzero & phi1)
			 | (OP==`ADC_zpx & T==`Tone & phi1)
			 | (OP==`ADC_zpx & T==`Ttwo & phi1)
			 | (OP==`ROR_zpx & T==`Tzero & phi1)
			 | (OP==`ROR_zpx & T==`Tone & phi1)
			 | (OP==`ROR_zpx & T==`Ttwo & phi1)
			 | (OP==`ROR_zpx & T==`Tfour & phi1)
			 | (OP==`ROR_zpx & T==`Tfive & phi1)
			 | (OP==`SEI & T==`Tone & phi1)
			 | (OP==`SEI & T==`Ttwo & phi1)
			 | (OP==`ADC_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ADC_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`ADC_aby & T==`Tone & phi1)
			 | (OP==`ADC_aby & T==`Ttwo & phi1)
			 | (OP==`ADC_aby & T==`Tthree & phi1)
			 | (OP==`ADC_aby & T==`Tfour & phi1)
			 | (OP==`ADC_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ADC_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`ADC_abx & T==`Tone & phi1)
			 | (OP==`ADC_abx & T==`Ttwo & phi1)
			 | (OP==`ADC_abx & T==`Tthree & phi1)
			 | (OP==`ADC_abx & T==`Tfour & phi1)
			 | (OP==`ROR_abx & T==`Tzero & phi1)
			 | (OP==`ROR_abx & T==`Tone & phi1)
			 | (OP==`ROR_abx & T==`Ttwo & phi1)
			 | (OP==`ROR_abx & T==`Tthree & phi1)
			 | (OP==`ROR_abx & T==`Tfour & phi1)
			 | (OP==`ROR_abx & T==`Tfive & phi1)
			 | (OP==`ROR_abx & T==`Tsix & phi1)
			 | (OP==`STA_izx & T==`Tzero & phi1)
			 | (OP==`STA_izx & T==`Tone & phi1)
			 | (OP==`STA_izx & T==`Ttwo & phi1)
			 | (OP==`STA_izx & T==`Tfive & phi1)
			 | (OP==`STY_zp & T==`Tone & phi1)
			 | (OP==`STY_zp & T==`Ttwo & phi1)
			 | (OP==`STA_zp & T==`Tone & phi1)
			 | (OP==`STA_zp & T==`Ttwo & phi1)
			 | (OP==`STX_zp & T==`Tone & phi1)
			 | (OP==`STX_zp & T==`Ttwo & phi1)
			 | (OP==`DEY & T==`Tone & phi1)
			 | (OP==`DEY & T==`Ttwo & phi1)
			 | (OP==`TXA & T==`Tone & phi1)
			 | (OP==`TXA & T==`Ttwo & phi1)
			 | (OP==`STY_abs & T==`Tzero & phi1)
			 | (OP==`STY_abs & T==`Tone & phi1)
			 | (OP==`STY_abs & T==`Ttwo & phi1)
			 | (OP==`STY_abs & T==`Tthree & phi1)
			 | (OP==`STA_abs & T==`Tzero & phi1)
			 | (OP==`STA_abs & T==`Tone & phi1)
			 | (OP==`STA_abs & T==`Ttwo & phi1)
			 | (OP==`STA_abs & T==`Tthree & phi1)
			 | (OP==`STX_abs & T==`Tzero & phi1)
			 | (OP==`STX_abs & T==`Tone & phi1)
			 | (OP==`STX_abs & T==`Ttwo & phi1)
			 | (OP==`STX_abs & T==`Tthree & phi1)
			 | (OP==`BCC_rel & T==`Ttwo & phi1)
			 | (OP==`BCC_rel & T==`T1BranchCross & phi1)
			 | (OP==`STA_izy & T==`Tzero & phi1)
			 | (OP==`STA_izy & T==`Tone & phi1)
			 | (OP==`STA_izy & T==`Ttwo & phi1)
			 | (OP==`STA_izy & T==`Tfour & phi1)
			 | (OP==`STA_izy & T==`Tfive & phi1)
			 | (OP==`STY_zpx & T==`Tzero & phi1)
			 | (OP==`STY_zpx & T==`Tone & phi1)
			 | (OP==`STY_zpx & T==`Ttwo & phi1)
			 | (OP==`STA_zpx & T==`Tzero & phi1)
			 | (OP==`STA_zpx & T==`Tone & phi1)
			 | (OP==`STA_zpx & T==`Ttwo & phi1)
			 | (OP==`STX_zpy & T==`Tzero & phi1)
			 | (OP==`STX_zpy & T==`Tone & phi1)
			 | (OP==`STX_zpy & T==`Ttwo & phi1)
			 | (OP==`TYA & T==`Tone & phi1)
			 | (OP==`TYA & T==`Ttwo & phi1)
			 | (OP==`STA_aby & T==`Tzero & phi1)
			 | (OP==`STA_aby & T==`Tone & phi1)
			 | (OP==`STA_aby & T==`Ttwo & phi1)
			 | (OP==`STA_aby & T==`Tthree & phi1)
			 | (OP==`STA_aby & T==`Tfour & phi1)
			 | (OP==`TXS & T==`Tone & phi1)
			 | (OP==`TXS & T==`Ttwo & phi1)
			 | (OP==`STA_abx & T==`Tzero & phi1)
			 | (OP==`STA_abx & T==`Tone & phi1)
			 | (OP==`STA_abx & T==`Ttwo & phi1)
			 | (OP==`STA_abx & T==`Tthree & phi1)
			 | (OP==`STA_abx & T==`Tfour & phi1)
			 | (OP==`LDY_imm & T==`Tone & phi1)
			 | (OP==`LDY_imm & T==`Ttwo & phi1)
			 | (OP==`LDA_izx & T==`Tzero & phi1)
			 | (OP==`LDA_izx & T==`Tone & phi1)
			 | (OP==`LDA_izx & T==`Ttwo & phi1)
			 | (OP==`LDA_izx & T==`Tfive & phi1)
			 | (OP==`LDX_imm & T==`Tone & phi1)
			 | (OP==`LDX_imm & T==`Ttwo & phi1)
			 | (OP==`LDY_zp & T==`Tone & phi1)
			 | (OP==`LDY_zp & T==`Ttwo & phi1)
			 | (OP==`LDA_zp & T==`Tone & phi1)
			 | (OP==`LDA_zp & T==`Ttwo & phi1)
			 | (OP==`LDX_zp & T==`Tone & phi1)
			 | (OP==`LDX_zp & T==`Ttwo & phi1)
			 | (OP==`TAY & T==`Tone & phi1)
			 | (OP==`TAY & T==`Ttwo & phi1)
			 | (OP==`LDA_imm & T==`Tone & phi1)
			 | (OP==`LDA_imm & T==`Ttwo & phi1)
			 | (OP==`TAX & T==`Tone & phi1)
			 | (OP==`TAX & T==`Ttwo & phi1)
			 | (OP==`LDY_abs & T==`Tzero & phi1)
			 | (OP==`LDY_abs & T==`Tone & phi1)
			 | (OP==`LDY_abs & T==`Ttwo & phi1)
			 | (OP==`LDY_abs & T==`Tthree & phi1)
			 | (OP==`LDA_abs & T==`Tzero & phi1)
			 | (OP==`LDA_abs & T==`Tone & phi1)
			 | (OP==`LDA_abs & T==`Ttwo & phi1)
			 | (OP==`LDA_abs & T==`Tthree & phi1)
			 | (OP==`LDX_abs & T==`Tzero & phi1)
			 | (OP==`LDX_abs & T==`Tone & phi1)
			 | (OP==`LDX_abs & T==`Ttwo & phi1)
			 | (OP==`LDX_abs & T==`Tthree & phi1)
			 | (OP==`BCS_rel & T==`Ttwo & phi1)
			 | (OP==`BCS_rel & T==`T1BranchCross & phi1)
			 | (OP==`LDA_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDA_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`LDA_izy & T==`Tone & phi1)
			 | (OP==`LDA_izy & T==`Ttwo & phi1)
			 | (OP==`LDA_izy & T==`Tfour & phi1)
			 | (OP==`LDA_izy & T==`Tfive & phi1)
			 | (OP==`LDY_zpx & T==`Tzero & phi1)
			 | (OP==`LDY_zpx & T==`Tone & phi1)
			 | (OP==`LDY_zpx & T==`Ttwo & phi1)
			 | (OP==`LDA_zpx & T==`Tzero & phi1)
			 | (OP==`LDA_zpx & T==`Tone & phi1)
			 | (OP==`LDA_zpx & T==`Ttwo & phi1)
			 | (OP==`LDX_zpy & T==`Tzero & phi1)
			 | (OP==`LDX_zpy & T==`Tone & phi1)
			 | (OP==`LDX_zpy & T==`Ttwo & phi1)
			 | (OP==`CLV & T==`Tone & phi1)
			 | (OP==`CLV & T==`Ttwo & phi1)
			 | (OP==`LDA_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDA_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`LDA_aby & T==`Tone & phi1)
			 | (OP==`LDA_aby & T==`Ttwo & phi1)
			 | (OP==`LDA_aby & T==`Tthree & phi1)
			 | (OP==`LDA_aby & T==`Tfour & phi1)
			 | (OP==`TSX & T==`Tone & phi1)
			 | (OP==`TSX & T==`Ttwo & phi1)
			 | (OP==`LDY_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDY_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`LDY_abx & T==`Tone & phi1)
			 | (OP==`LDY_abx & T==`Ttwo & phi1)
			 | (OP==`LDY_abx & T==`Tthree & phi1)
			 | (OP==`LDY_abx & T==`Tfour & phi1)
			 | (OP==`LDA_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDA_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`LDA_abx & T==`Tone & phi1)
			 | (OP==`LDA_abx & T==`Ttwo & phi1)
			 | (OP==`LDA_abx & T==`Tthree & phi1)
			 | (OP==`LDA_abx & T==`Tfour & phi1)
			 | (OP==`LDX_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDX_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`LDX_aby & T==`Tone & phi1)
			 | (OP==`LDX_aby & T==`Ttwo & phi1)
			 | (OP==`LDX_aby & T==`Tthree & phi1)
			 | (OP==`LDX_aby & T==`Tfour & phi1)
			 | (OP==`CPY_imm & T==`Ttwo & phi1)
			 | (OP==`CMP_izx & T==`Tzero & phi1)
			 | (OP==`CMP_izx & T==`Ttwo & phi1)
			 | (OP==`CMP_izx & T==`Tfive & phi1)
			 | (OP==`CPY_zp & T==`Ttwo & phi1)
			 | (OP==`CMP_zp & T==`Ttwo & phi1)
			 | (OP==`DEC_zp & T==`Tzero & phi1)
			 | (OP==`DEC_zp & T==`Tone & phi1)
			 | (OP==`DEC_zp & T==`Ttwo & phi1)
			 | (OP==`DEC_zp & T==`Tfour & phi1)
			 | (OP==`INY & T==`Ttwo & phi1)
			 | (OP==`CMP_imm & T==`Ttwo & phi1)
			 | (OP==`DEX & T==`Tone & phi1)
			 | (OP==`DEX & T==`Ttwo & phi1)
			 | (OP==`CPY_abs & T==`Tzero & phi1)
			 | (OP==`CPY_abs & T==`Ttwo & phi1)
			 | (OP==`CPY_abs & T==`Tthree & phi1)
			 | (OP==`CMP_abs & T==`Tzero & phi1)
			 | (OP==`CMP_abs & T==`Ttwo & phi1)
			 | (OP==`CMP_abs & T==`Tthree & phi1)
			 | (OP==`DEC_abs & T==`Tzero & phi1)
			 | (OP==`DEC_abs & T==`Tone & phi1)
			 | (OP==`DEC_abs & T==`Ttwo & phi1)
			 | (OP==`DEC_abs & T==`Tthree & phi1)
			 | (OP==`DEC_abs & T==`Tfour & phi1)
			 | (OP==`DEC_abs & T==`Tfive & phi1)
			 | (OP==`BNE_rel & T==`Ttwo & phi1)
			 | (OP==`BNE_rel & T==`T1BranchCross & phi1)
			 | (OP==`CMP_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`CMP_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`CMP_izy & T==`Ttwo & phi1)
			 | (OP==`CMP_izy & T==`Tfour & phi1)
			 | (OP==`CMP_izy & T==`Tfive & phi1)
			 | (OP==`CMP_zpx & T==`Tzero & phi1)
			 | (OP==`CMP_zpx & T==`Ttwo & phi1)
			 | (OP==`DEC_zpx & T==`Tzero & phi1)
			 | (OP==`DEC_zpx & T==`Tone & phi1)
			 | (OP==`DEC_zpx & T==`Ttwo & phi1)
			 | (OP==`DEC_zpx & T==`Tfour & phi1)
			 | (OP==`DEC_zpx & T==`Tfive & phi1)
			 | (OP==`CLD & T==`Tone & phi1)
			 | (OP==`CLD & T==`Ttwo & phi1)
			 | (OP==`CMP_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`CMP_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`CMP_aby & T==`Ttwo & phi1)
			 | (OP==`CMP_aby & T==`Tthree & phi1)
			 | (OP==`CMP_aby & T==`Tfour & phi1)
			 | (OP==`CMP_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`CMP_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`CMP_abx & T==`Ttwo & phi1)
			 | (OP==`CMP_abx & T==`Tthree & phi1)
			 | (OP==`CMP_abx & T==`Tfour & phi1)
			 | (OP==`DEC_abx & T==`Tzero & phi1)
			 | (OP==`DEC_abx & T==`Tone & phi1)
			 | (OP==`DEC_abx & T==`Ttwo & phi1)
			 | (OP==`DEC_abx & T==`Tthree & phi1)
			 | (OP==`DEC_abx & T==`Tfour & phi1)
			 | (OP==`DEC_abx & T==`Tfive & phi1)
			 | (OP==`DEC_abx & T==`Tsix & phi1)
			 | (OP==`CPX_imm & T==`Ttwo & phi1)
			 | (OP==`SBC_izx & T==`Tzero & phi1)
			 | (OP==`SBC_izx & T==`Ttwo & phi1)
			 | (OP==`SBC_izx & T==`Tfive & phi1)
			 | (OP==`CPX_zp & T==`Ttwo & phi1)
			 | (OP==`SBC_zp & T==`Ttwo & phi1)
			 | (OP==`INC_zp & T==`Tzero & phi1)
			 | (OP==`INC_zp & T==`Tone & phi1)
			 | (OP==`INC_zp & T==`Ttwo & phi1)
			 | (OP==`INC_zp & T==`Tfour & phi1)
			 | (OP==`INX & T==`Ttwo & phi1)
			 | (OP==`SBC_imm & T==`Ttwo & phi1)
			 | (OP==`NOP & T==`Tone & phi1)
			 | (OP==`NOP & T==`Ttwo & phi1)
			 | (OP==`CPX_abs & T==`Tzero & phi1)
			 | (OP==`CPX_abs & T==`Ttwo & phi1)
			 | (OP==`CPX_abs & T==`Tthree & phi1)
			 | (OP==`SBC_abs & T==`Tzero & phi1)
			 | (OP==`SBC_abs & T==`Ttwo & phi1)
			 | (OP==`SBC_abs & T==`Tthree & phi1)
			 | (OP==`INC_abs & T==`Tzero & phi1)
			 | (OP==`INC_abs & T==`Tone & phi1)
			 | (OP==`INC_abs & T==`Ttwo & phi1)
			 | (OP==`INC_abs & T==`Tthree & phi1)
			 | (OP==`INC_abs & T==`Tfour & phi1)
			 | (OP==`INC_abs & T==`Tfive & phi1)
			 | (OP==`BEQ_rel & T==`Ttwo & phi1)
			 | (OP==`BEQ_rel & T==`T1BranchCross & phi1)
			 | (OP==`SBC_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`SBC_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`SBC_izy & T==`Ttwo & phi1)
			 | (OP==`SBC_izy & T==`Tfour & phi1)
			 | (OP==`SBC_izy & T==`Tfive & phi1)
			 | (OP==`SBC_zpx & T==`Tzero & phi1)
			 | (OP==`SBC_zpx & T==`Ttwo & phi1)
			 | (OP==`INC_zpx & T==`Tzero & phi1)
			 | (OP==`INC_zpx & T==`Tone & phi1)
			 | (OP==`INC_zpx & T==`Ttwo & phi1)
			 | (OP==`INC_zpx & T==`Tfour & phi1)
			 | (OP==`INC_zpx & T==`Tfive & phi1)
			 | (OP==`SED & T==`Tone & phi1)
			 | (OP==`SED & T==`Ttwo & phi1)
			 | (OP==`SBC_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`SBC_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`SBC_aby & T==`Ttwo & phi1)
			 | (OP==`SBC_aby & T==`Tthree & phi1)
			 | (OP==`SBC_aby & T==`Tfour & phi1)
			 | (OP==`SBC_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`SBC_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`SBC_abx & T==`Ttwo & phi1)
			 | (OP==`SBC_abx & T==`Tthree & phi1)
			 | (OP==`SBC_abx & T==`Tfour & phi1)
			 | (OP==`INC_abx & T==`Tzero & phi1)
			 | (OP==`INC_abx & T==`Tone & phi1)
			 | (OP==`INC_abx & T==`Ttwo & phi1)
			 | (OP==`INC_abx & T==`Tthree & phi1)
			 | (OP==`INC_abx & T==`Tfour & phi1)
			 | (OP==`INC_abx & T==`Tfive & phi1)
			 | (OP==`INC_abx & T==`Tsix & phi1)
			;

assign control[`ADL_ADD] = (OP==`BRK & T==`Tthree & phi1)
			 | (OP==`BRK & T==`Tfour & phi1)
			 | (OP==`BRK & T==`Tfive & phi1)
			 | (OP==`ORA_izx & T==`Tthree & phi1)
			 | (OP==`ORA_izx & T==`Tfour & phi1)
			 | (OP==`ORA_zp & T==`Tzero & phi1)
			 | (OP==`ASL_zp & T==`Tthree & phi1)
			 | (OP==`PHP & T==`Tzero & phi1)
			 | (OP==`BPL_rel & T==`Tthree & phi1)
			 | (OP==`BPL_rel & T==`T1NoBranch & phi1)
			 | (OP==`ORA_izy & T==`Tthree & phi1)
			 | (OP==`ORA_zpx & T==`Tthree & phi1)
			 | (OP==`ASL_zpx & T==`Tthree & phi1)
			 | (OP==`JSR_abs & T==`Tthree & phi1)
			 | (OP==`JSR_abs & T==`Tfour & phi1)
			 | (OP==`JSR_abs & T==`Tfive & phi1)
			 | (OP==`AND_izx & T==`Tthree & phi1)
			 | (OP==`AND_izx & T==`Tfour & phi1)
			 | (OP==`BIT_zp & T==`Tzero & phi1)
			 | (OP==`AND_zp & T==`Tzero & phi1)
			 | (OP==`ROL_zp & T==`Tthree & phi1)
			 | (OP==`PLP & T==`Tzero & phi1)
			 | (OP==`PLP & T==`Tthree & phi1)
			 | (OP==`BIT_abs & T==`Tzero & phi1)
			 | (OP==`BMI_rel & T==`Tthree & phi1)
			 | (OP==`BMI_rel & T==`T1NoBranch & phi1)
			 | (OP==`AND_izy & T==`Tthree & phi1)
			 | (OP==`AND_zpx & T==`Tthree & phi1)
			 | (OP==`ROL_zpx & T==`Tthree & phi1)
			 | (OP==`RTI & T==`Tthree & phi1)
			 | (OP==`RTI & T==`Tfour & phi1)
			 | (OP==`RTI & T==`Tfive & phi1)
			 | (OP==`EOR_izx & T==`Tthree & phi1)
			 | (OP==`EOR_izx & T==`Tfour & phi1)
			 | (OP==`EOR_zp & T==`Tzero & phi1)
			 | (OP==`LSR_zp & T==`Tthree & phi1)
			 | (OP==`PHA & T==`Tzero & phi1)
			 | (OP==`BVC_rel & T==`Tthree & phi1)
			 | (OP==`BVC_rel & T==`T1NoBranch & phi1)
			 | (OP==`EOR_izy & T==`Tthree & phi1)
			 | (OP==`EOR_zpx & T==`Tthree & phi1)
			 | (OP==`LSR_zpx & T==`Tthree & phi1)
			 | (OP==`RTS & T==`Tthree & phi1)
			 | (OP==`RTS & T==`Tfour & phi1)
			 | (OP==`ADC_izx & T==`Tthree & phi1)
			 | (OP==`ADC_izx & T==`Tfour & phi1)
			 | (OP==`ADC_zp & T==`Tzero & phi1)
			 | (OP==`ROR_zp & T==`Tthree & phi1)
			 | (OP==`PLA & T==`Tzero & phi1)
			 | (OP==`PLA & T==`Tthree & phi1)
			 | (OP==`JMP_zp & T==`Tfour & phi1)
			 | (OP==`BVS_rel & T==`Tthree & phi1)
			 | (OP==`BVS_rel & T==`T1NoBranch & phi1)
			 | (OP==`ADC_izy & T==`Tthree & phi1)
			 | (OP==`ADC_zpx & T==`Tthree & phi1)
			 | (OP==`ROR_zpx & T==`Tthree & phi1)
			 | (OP==`STA_izx & T==`Tthree & phi1)
			 | (OP==`STA_izx & T==`Tfour & phi1)
			 | (OP==`STY_zp & T==`Tzero & phi1)
			 | (OP==`STA_zp & T==`Tzero & phi1)
			 | (OP==`STX_zp & T==`Tzero & phi1)
			 | (OP==`BCC_rel & T==`Tthree & phi1)
			 | (OP==`BCC_rel & T==`T1NoBranch & phi1)
			 | (OP==`STA_izy & T==`Tthree & phi1)
			 | (OP==`STY_zpx & T==`Tthree & phi1)
			 | (OP==`STA_zpx & T==`Tthree & phi1)
			 | (OP==`STX_zpy & T==`Tthree & phi1)
			 | (OP==`LDA_izx & T==`Tthree & phi1)
			 | (OP==`LDA_izx & T==`Tfour & phi1)
			 | (OP==`LDY_zp & T==`Tzero & phi1)
			 | (OP==`LDA_zp & T==`Tzero & phi1)
			 | (OP==`LDX_zp & T==`Tzero & phi1)
			 | (OP==`BCS_rel & T==`Tthree & phi1)
			 | (OP==`BCS_rel & T==`T1NoBranch & phi1)
			 | (OP==`LDA_izy & T==`Tthree & phi1)
			 | (OP==`LDY_zpx & T==`Tthree & phi1)
			 | (OP==`LDA_zpx & T==`Tthree & phi1)
			 | (OP==`LDX_zpy & T==`Tthree & phi1)
			 | (OP==`CMP_izx & T==`Tthree & phi1)
			 | (OP==`CMP_izx & T==`Tfour & phi1)
			 | (OP==`CPY_zp & T==`Tzero & phi1)
			 | (OP==`CMP_zp & T==`Tzero & phi1)
			 | (OP==`DEC_zp & T==`Tthree & phi1)
			 | (OP==`BNE_rel & T==`Tthree & phi1)
			 | (OP==`BNE_rel & T==`T1NoBranch & phi1)
			 | (OP==`CMP_izy & T==`Tthree & phi1)
			 | (OP==`CMP_zpx & T==`Tthree & phi1)
			 | (OP==`DEC_zpx & T==`Tthree & phi1)
			 | (OP==`SBC_izx & T==`Tthree & phi1)
			 | (OP==`SBC_izx & T==`Tfour & phi1)
			 | (OP==`CPX_zp & T==`Tzero & phi1)
			 | (OP==`SBC_zp & T==`Tzero & phi1)
			 | (OP==`INC_zp & T==`Tthree & phi1)
			 | (OP==`BEQ_rel & T==`Tthree & phi1)
			 | (OP==`BEQ_rel & T==`T1NoBranch & phi1)
			 | (OP==`SBC_izy & T==`Tthree & phi1)
			 | (OP==`SBC_zpx & T==`Tthree & phi1)
			 | (OP==`INC_zpx & T==`Tthree & phi1)
			;

assign control[`I_ADDC] = (OP==`ORA_izx & T==`Tfour)
			 | (OP==`ORA_izx & T==`Tfour & phi1)
			 | (OP==`ORA_izx & T==`Tfour & phi2)
			 | (OP==`BPL_rel & T==`Tzero & phi1)
			 | (OP==`BPL_rel & T==`Tzero & phi2)
			 | (OP==`BPL_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BPL_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`ORA_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ORA_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`ORA_izy & T==`Tthree & phi1)
			 | (OP==`ORA_izy & T==`Tthree & phi2)
			 | (OP==`ORA_izy & T==`Tfive & phi1)
			 | (OP==`ORA_izy & T==`Tfive & phi2)
			 | (OP==`ORA_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ORA_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`ORA_aby & T==`Tfour & phi1)
			 | (OP==`ORA_aby & T==`Tfour & phi2)
			 | (OP==`ORA_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ORA_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`ORA_abx & T==`Tfour & phi1)
			 | (OP==`ORA_abx & T==`Tfour & phi2)
			 | (OP==`ASL_abx & T==`Tfour & phi1)
			 | (OP==`ASL_abx & T==`Tfour & phi2)
			 | (OP==`AND_izx & T==`Tfour & phi1)
			 | (OP==`AND_izx & T==`Tfour & phi2)
			 | (OP==`ROL_zp & T==`Tfour & phi1 & statusC)
			 | (OP==`ROL_zp & T==`Tfour & phi2 & statusC)
			 | (OP==`PLP & T==`Tzero & phi1)
			 | (OP==`PLP & T==`Tzero & phi2)
			 | (OP==`PLP & T==`Tthree & phi1)
			 | (OP==`PLP & T==`Tthree & phi2)
			 | (OP==`ROL & T==`Tone & phi1 & statusC)
			 | (OP==`ROL & T==`Tone & phi2 & statusC)
			 | (OP==`ROL_abs & T==`Tfive & phi1 & statusC)
			 | (OP==`ROL_abs & T==`Tfive & phi2 & statusC)
			 | (OP==`BMI_rel & T==`Tzero & phi1)
			 | (OP==`BMI_rel & T==`Tzero & phi2)
			 | (OP==`BMI_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BMI_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`AND_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`AND_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`AND_izy & T==`Tthree & phi1)
			 | (OP==`AND_izy & T==`Tthree & phi2)
			 | (OP==`AND_izy & T==`Tfive & phi1)
			 | (OP==`AND_izy & T==`Tfive & phi2)
			 | (OP==`ROL_zpx & T==`Tfive & phi1 & statusC)
			 | (OP==`ROL_zpx & T==`Tfive & phi2 & statusC)
			 | (OP==`AND_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`AND_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`AND_aby & T==`Tfour & phi1)
			 | (OP==`AND_aby & T==`Tfour & phi2)
			 | (OP==`AND_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`AND_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`AND_abx & T==`Tfour & phi1)
			 | (OP==`AND_abx & T==`Tfour & phi2)
			 | (OP==`ROL_abx & T==`Tfour & phi1)
			 | (OP==`ROL_abx & T==`Tfour & phi2)
			 | (OP==`ROL_abx & T==`Tsix & phi1 & statusC)
			 | (OP==`ROL_abx & T==`Tsix & phi2 & statusC)
			 | (OP==`RTI & T==`Tthree & phi1)
			 | (OP==`RTI & T==`Tthree & phi2)
			 | (OP==`RTI & T==`Tfour & phi1)
			 | (OP==`RTI & T==`Tfour & phi2)
			 | (OP==`RTI & T==`Tfive & phi1)
			 | (OP==`RTI & T==`Tfive & phi2)
			 | (OP==`EOR_izx & T==`Tfour & phi1)
			 | (OP==`EOR_izx & T==`Tfour & phi2)
			 | (OP==`BVC_rel & T==`Tzero & phi1)
			 | (OP==`BVC_rel & T==`Tzero & phi2)
			 | (OP==`BVC_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BVC_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`EOR_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`EOR_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`EOR_izy & T==`Tthree & phi1)
			 | (OP==`EOR_izy & T==`Tthree & phi2)
			 | (OP==`EOR_izy & T==`Tfive & phi1)
			 | (OP==`EOR_izy & T==`Tfive & phi2)
			 | (OP==`EOR_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`EOR_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`EOR_aby & T==`Tfour & phi1)
			 | (OP==`EOR_aby & T==`Tfour & phi2)
			 | (OP==`EOR_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`EOR_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`EOR_abx & T==`Tfour & phi1)
			 | (OP==`EOR_abx & T==`Tfour & phi2)
			 | (OP==`LSR_abx & T==`Tfour & phi1)
			 | (OP==`LSR_abx & T==`Tfour & phi2)
			 | (OP==`RTS & T==`Tthree & phi1)
			 | (OP==`RTS & T==`Tthree & phi2)
			 | (OP==`RTS & T==`Tfour & phi1)
			 | (OP==`RTS & T==`Tfour & phi2)
			 | (OP==`ADC_izx & T==`Tone & phi1 & statusC)
			 | (OP==`ADC_izx & T==`Tone & phi2 & statusC)
			 | (OP==`ADC_izx & T==`Tfour & phi1)
			 | (OP==`ADC_izx & T==`Tfour & phi2)
			 | (OP==`ADC_zp & T==`Tone & phi1 & statusC)
			 | (OP==`ADC_zp & T==`Tone & phi2 & statusC)
			 | (OP==`ROR_zp & T==`Tfour & phi1 & statusC)
			 | (OP==`ROR_zp & T==`Tfour & phi2 & statusC)
			 | (OP==`PLA & T==`Tzero & phi1)
			 | (OP==`PLA & T==`Tzero & phi2)
			 | (OP==`PLA & T==`Tthree & phi1)
			 | (OP==`PLA & T==`Tthree & phi2)
			 | (OP==`ADC_imm & T==`Tone & phi1 & statusC)
			 | (OP==`ADC_imm & T==`Tone & phi2 & statusC)
			 | (OP==`ROR & T==`Tone & phi1 & statusC)
			 | (OP==`ROR & T==`Tone & phi2 & statusC)
			 | (OP==`JMP_zp & T==`Tfour & phi1)
			 | (OP==`JMP_zp & T==`Tfour & phi2)
			 | (OP==`ADC_abs & T==`Tone & phi1 & statusC)
			 | (OP==`ADC_abs & T==`Tone & phi2 & statusC)
			 | (OP==`ROR_abs & T==`Tfive & phi1 & statusC)
			 | (OP==`ROR_abs & T==`Tfive & phi2 & statusC)
			 | (OP==`BVS_rel & T==`Tzero & phi1)
			 | (OP==`BVS_rel & T==`Tzero & phi2)
			 | (OP==`BVS_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BVS_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`ADC_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ADC_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`ADC_izy & T==`Tone & phi1 & statusC)
			 | (OP==`ADC_izy & T==`Tone & phi2 & statusC)
			 | (OP==`ADC_izy & T==`Tthree & phi1)
			 | (OP==`ADC_izy & T==`Tthree & phi2)
			 | (OP==`ADC_izy & T==`Tfive & phi1)
			 | (OP==`ADC_izy & T==`Tfive & phi2)
			 | (OP==`ADC_zpx & T==`Tone & phi1 & statusC)
			 | (OP==`ADC_zpx & T==`Tone & phi2 & statusC)
			 | (OP==`ROR_zpx & T==`Tfive & phi1 & statusC)
			 | (OP==`ROR_zpx & T==`Tfive & phi2 & statusC)
			 | (OP==`ADC_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ADC_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`ADC_aby & T==`Tone & phi1 & statusC)
			 | (OP==`ADC_aby & T==`Tone & phi2 & statusC)
			 | (OP==`ADC_aby & T==`Tfour & phi2)
			 | (OP==`ADC_abx & T==`Tone & phi1 & statusC)
			 | (OP==`ADC_abx & T==`Tone & phi2 & statusC)
			 | (OP==`ROR_abx & T==`Tfour & phi1)
			 | (OP==`ROR_abx & T==`Tfour & phi2)
			 | (OP==`ROR_abx & T==`Tsix & phi1 & statusC)
			 | (OP==`ROR_abx & T==`Tsix & phi2 & statusC)
			 | (OP==`STA_izx & T==`Tfour & phi1)
			 | (OP==`STA_izx & T==`Tfour & phi2)
			 | (OP==`BCC_rel & T==`Tzero & phi1)
			 | (OP==`BCC_rel & T==`Tzero & phi2)
			 | (OP==`BCC_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BCC_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`STA_izy & T==`Tthree & phi1)
			 | (OP==`STA_izy & T==`Tthree & phi2)
			 | (OP==`STA_izy & T==`Tfive & phi1)
			 | (OP==`STA_izy & T==`Tfive & phi2)
			 | (OP==`STA_aby & T==`Tfour & phi1)
			 | (OP==`STA_aby & T==`Tfour & phi2)
			 | (OP==`STA_abx & T==`Tfour & phi1)
			 | (OP==`STA_abx & T==`Tfour & phi2)
			 | (OP==`LDA_izx & T==`Tfour & phi1)
			 | (OP==`LDA_izx & T==`Tfour & phi2)
			 | (OP==`BCS_rel & T==`Tzero & phi1)
			 | (OP==`BCS_rel & T==`Tzero & phi2)
			 | (OP==`BCS_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BCS_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`LDA_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDA_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`LDA_izy & T==`Tthree & phi1)
			 | (OP==`LDA_izy & T==`Tthree & phi2)
			 | (OP==`LDA_izy & T==`Tfive & phi1)
			 | (OP==`LDA_izy & T==`Tfive & phi2)
			 | (OP==`LDA_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDA_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`LDA_aby & T==`Tfour & phi1)
			 | (OP==`LDA_aby & T==`Tfour & phi2)
			 | (OP==`LDY_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDY_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`LDY_abx & T==`Tfour & phi1)
			 | (OP==`LDY_abx & T==`Tfour & phi2)
			 | (OP==`LDA_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDA_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`LDA_abx & T==`Tfour & phi1)
			 | (OP==`LDA_abx & T==`Tfour & phi2)
			 | (OP==`LDX_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDX_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`LDX_aby & T==`Tfour & phi1)
			 | (OP==`LDX_aby & T==`Tfour & phi2)
			 | (OP==`CPY_imm & T==`Tone & phi1)
			 | (OP==`CPY_imm & T==`Tone & phi2)
			 | (OP==`CMP_izx & T==`Tfour & phi1)
			 | (OP==`CMP_izx & T==`Tfour & phi2)
			 | (OP==`CPY_zp & T==`Tone & phi1)
			 | (OP==`CPY_zp & T==`Tone & phi2)
			 | (OP==`CMP_zp & T==`Tone & phi1)
			 | (OP==`CMP_zp & T==`Tone & phi1)
			 | (OP==`CMP_zp & T==`Tone & phi2)
			 | (OP==`CMP_zp & T==`Tone & phi2)
			 | (OP==`INY & T==`Tone & phi1)
			 | (OP==`INY & T==`Tone & phi2)
			 | (OP==`CMP_imm & T==`Tone & phi1)
			 | (OP==`CMP_imm & T==`Tone & phi2)
			 | (OP==`CPY_abs & T==`Tone & phi1)
			 | (OP==`CPY_abs & T==`Tone & phi2)
			 | (OP==`CMP_abs & T==`Tone & phi1)
			 | (OP==`CMP_abs & T==`Tone & phi2)
			 | (OP==`BNE_rel & T==`Tzero & phi1)
			 | (OP==`BNE_rel & T==`Tzero & phi2)
			 | (OP==`BNE_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BNE_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`CMP_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`CMP_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`CMP_izy & T==`Tone & phi1)
			 | (OP==`CMP_izy & T==`Tone & phi2)
			 | (OP==`CMP_izy & T==`Tthree & phi1)
			 | (OP==`CMP_izy & T==`Tthree & phi2)
			 | (OP==`CMP_izy & T==`Tfive & phi1)
			 | (OP==`CMP_izy & T==`Tfive & phi2)
			 | (OP==`CMP_zpx & T==`Tone & phi1)
			 | (OP==`CMP_zpx & T==`Tone & phi2)
			 | (OP==`CMP_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`CMP_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`CMP_aby & T==`Tone & phi1)
			 | (OP==`CMP_aby & T==`Tone & phi2)
			 | (OP==`CMP_aby & T==`Tfour & phi1)
			 | (OP==`CMP_aby & T==`Tfour & phi2)
			 | (OP==`CMP_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`CMP_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`CMP_abx & T==`Tone & phi1)
			 | (OP==`CMP_abx & T==`Tone & phi2)
			 | (OP==`CMP_abx & T==`Tfour & phi1)
			 | (OP==`CMP_abx & T==`Tfour & phi2)
			 | (OP==`DEC_abx & T==`Tfour & phi1)
			 | (OP==`DEC_abx & T==`Tfour & phi2)
			 | (OP==`CPX_imm & T==`Tone & phi1)
			 | (OP==`CPX_imm & T==`Tone & phi2)
			 | (OP==`SBC_izx & T==`Tone & phi1 & statusC)
			 | (OP==`SBC_izx & T==`Tone & phi2 & statusC)
			 | (OP==`SBC_izx & T==`Tfour & phi1)
			 | (OP==`SBC_izx & T==`Tfour & phi2)
			 | (OP==`CPX_zp & T==`Tone & phi1)
			 | (OP==`CPX_zp & T==`Tone & phi2)
			 | (OP==`SBC_zp & T==`Tone & phi1 & statusC)
			 | (OP==`SBC_zp & T==`Tone & phi2 & statusC)
			 | (OP==`INC_zp & T==`Tfour & phi1)
			 | (OP==`INC_zp & T==`Tfour & phi2)
			 | (OP==`INX & T==`Tone & phi1)
			 | (OP==`INX & T==`Tone & phi2)
			 | (OP==`SBC_imm & T==`Tone & phi1 & statusC)
			 | (OP==`SBC_imm & T==`Tone & phi2 & statusC)
			 | (OP==`CPX_abs & T==`Tone & phi1)
			 | (OP==`CPX_abs & T==`Tone & phi2)
			 | (OP==`SBC_abs & T==`Tone & phi1 & statusC)
			 | (OP==`SBC_abs & T==`Tone & phi2 & statusC)
			 | (OP==`INC_abs & T==`Tfive & phi1)
			 | (OP==`INC_abs & T==`Tfive & phi2)
			 | (OP==`BEQ_rel & T==`Tzero & phi1)
			 | (OP==`BEQ_rel & T==`Tzero & phi2)
			 | (OP==`BEQ_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BEQ_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`SBC_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`SBC_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`SBC_izy & T==`Tone & phi1 & statusC)
			 | (OP==`SBC_izy & T==`Tone & phi2 & statusC)
			 | (OP==`SBC_izy & T==`Tthree & phi1)
			 | (OP==`SBC_izy & T==`Tthree & phi2)
			 | (OP==`SBC_izy & T==`Tfive & phi1)
			 | (OP==`SBC_izy & T==`Tfive & phi2)
			 | (OP==`SBC_zpx & T==`Tone & phi1 & statusC)
			 | (OP==`SBC_zpx & T==`Tone & phi2 & statusC)
			 | (OP==`INC_zpx & T==`Tfive & phi1)
			 | (OP==`INC_zpx & T==`Tfive & phi2)
			 | (OP==`SBC_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`SBC_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`SBC_aby & T==`Tone & phi1 & statusC)
			 | (OP==`SBC_aby & T==`Tone & phi2 & statusC)
			 | (OP==`SBC_aby & T==`Tfour & phi1)
			 | (OP==`SBC_aby & T==`Tfour & phi2)
			 | (OP==`SBC_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`SBC_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`SBC_abx & T==`Tone & phi1 & statusC)
			 | (OP==`SBC_abx & T==`Tone & phi2 & statusC)
			 | (OP==`SBC_abx & T==`Tfour & phi1)
			 | (OP==`SBC_abx & T==`Tfour & phi2)
			 | (OP==`INC_abx & T==`Tfour & phi1)
			 | (OP==`INC_abx & T==`Tfour & phi2)
			 | (OP==`INC_abx & T==`Tsix & phi1)
			 | (OP==`INC_abx & T==`Tsix & phi2)
			;

assign control[`nDAA] = (OP==`BRK & T==`Tzero & phi1)
			 | (OP==`BRK & T==`Tzero & phi2)
			 | (OP==`BRK & T==`Tone & phi1)
			 | (OP==`BRK & T==`Tone & phi2)
			 | (OP==`BRK & T==`Ttwo & phi1)
			 | (OP==`BRK & T==`Ttwo & phi2)
			 | (OP==`BRK & T==`Tthree & phi1)
			 | (OP==`BRK & T==`Tthree & phi2)
			 | (OP==`BRK & T==`Tfour & phi1)
			 | (OP==`BRK & T==`Tfour & phi2)
			 | (OP==`BRK & T==`Tfive & phi1)
			 | (OP==`BRK & T==`Tfive & phi2)
			 | (OP==`BRK & T==`Tsix & phi1)
			 | (OP==`BRK & T==`Tsix & phi2)
			 | (OP==`ORA_izx & T==`Tzero & phi1)
			 | (OP==`ORA_izx & T==`Tzero & phi2)
			 | (OP==`ORA_izx & T==`Tone & phi1)
			 | (OP==`ORA_izx & T==`Tone & phi2)
			 | (OP==`ORA_izx & T==`Ttwo & phi1)
			 | (OP==`ORA_izx & T==`Ttwo & phi2)
			 | (OP==`ORA_izx & T==`Tthree & phi1)
			 | (OP==`ORA_izx & T==`Tthree & phi2)
			 | (OP==`ORA_izx & T==`Tfour & phi1)
			 | (OP==`ORA_izx & T==`Tfour & phi2)
			 | (OP==`ORA_izx & T==`Tfive & phi1)
			 | (OP==`ORA_izx & T==`Tfive & phi2)
			 | (OP==`ORA_zp & T==`Tzero & phi1)
			 | (OP==`ORA_zp & T==`Tzero & phi2)
			 | (OP==`ORA_zp & T==`Tone & phi1)
			 | (OP==`ORA_zp & T==`Tone & phi2)
			 | (OP==`ORA_zp & T==`Ttwo & phi1)
			 | (OP==`ORA_zp & T==`Ttwo & phi2)
			 | (OP==`ASL_zp & T==`Tzero & phi1)
			 | (OP==`ASL_zp & T==`Tzero & phi2)
			 | (OP==`ASL_zp & T==`Tone & phi1)
			 | (OP==`ASL_zp & T==`Tone & phi2)
			 | (OP==`ASL_zp & T==`Ttwo & phi1)
			 | (OP==`ASL_zp & T==`Ttwo & phi2)
			 | (OP==`ASL_zp & T==`Tthree & phi1)
			 | (OP==`ASL_zp & T==`Tthree & phi2)
			 | (OP==`ASL_zp & T==`Tfour & phi1)
			 | (OP==`ASL_zp & T==`Tfour & phi2)
			 | (OP==`PHP & T==`Tzero & phi1)
			 | (OP==`PHP & T==`Tzero & phi2)
			 | (OP==`PHP & T==`Tone & phi1)
			 | (OP==`PHP & T==`Tone & phi2)
			 | (OP==`PHP & T==`Ttwo & phi1)
			 | (OP==`PHP & T==`Ttwo & phi2)
			 | (OP==`ORA_imm & T==`Tone & phi1)
			 | (OP==`ORA_imm & T==`Tone & phi2)
			 | (OP==`ORA_imm & T==`Ttwo & phi1)
			 | (OP==`ORA_imm & T==`Ttwo & phi2)
			 | (OP==`ASL & T==`Tone & phi1)
			 | (OP==`ASL & T==`Tone & phi2)
			 | (OP==`ASL & T==`Ttwo & phi1)
			 | (OP==`ASL & T==`Ttwo & phi2)
			 | (OP==`ORA_abs & T==`Tzero & phi1)
			 | (OP==`ORA_abs & T==`Tzero & phi2)
			 | (OP==`ORA_abs & T==`Tone & phi1)
			 | (OP==`ORA_abs & T==`Tone & phi2)
			 | (OP==`ORA_abs & T==`Ttwo & phi1)
			 | (OP==`ORA_abs & T==`Ttwo & phi2)
			 | (OP==`ORA_abs & T==`Tthree & phi1)
			 | (OP==`ORA_abs & T==`Tthree & phi2)
			 | (OP==`ASL_abs & T==`Tzero & phi1)
			 | (OP==`ASL_abs & T==`Tzero & phi2)
			 | (OP==`ASL_abs & T==`Tone & phi1)
			 | (OP==`ASL_abs & T==`Tone & phi2)
			 | (OP==`ASL_abs & T==`Ttwo & phi1)
			 | (OP==`ASL_abs & T==`Ttwo & phi2)
			 | (OP==`ASL_abs & T==`Tthree & phi1)
			 | (OP==`ASL_abs & T==`Tthree & phi2)
			 | (OP==`ASL_abs & T==`Tfour & phi1)
			 | (OP==`ASL_abs & T==`Tfour & phi2)
			 | (OP==`ASL_abs & T==`Tfive & phi1)
			 | (OP==`ASL_abs & T==`Tfive & phi2)
			 | (OP==`BPL_rel & T==`Tzero & phi1)
			 | (OP==`BPL_rel & T==`Tzero & phi2)
			 | (OP==`BPL_rel & T==`Ttwo & phi1)
			 | (OP==`BPL_rel & T==`Ttwo & phi2)
			 | (OP==`BPL_rel & T==`Tthree & phi1)
			 | (OP==`BPL_rel & T==`Tthree & phi2)
			 | (OP==`BPL_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BPL_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BPL_rel & T==`T1BranchCross & phi1)
			 | (OP==`BPL_rel & T==`T1BranchCross & phi2)
			 | (OP==`BPL_rel & T==`T1NoBranch & phi1)
			 | (OP==`BPL_rel & T==`T1NoBranch & phi2)
			 | (OP==`ORA_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`ORA_izy & T==`TzeroCrossPg & phi2)
			 | (OP==`ORA_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ORA_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`ORA_izy & T==`Tone & phi1)
			 | (OP==`ORA_izy & T==`Tone & phi2)
			 | (OP==`ORA_izy & T==`Ttwo & phi1)
			 | (OP==`ORA_izy & T==`Ttwo & phi2)
			 | (OP==`ORA_izy & T==`Tthree & phi1)
			 | (OP==`ORA_izy & T==`Tthree & phi2)
			 | (OP==`ORA_izy & T==`Tfour & phi1)
			 | (OP==`ORA_izy & T==`Tfour & phi2)
			 | (OP==`ORA_izy & T==`Tfive & phi1)
			 | (OP==`ORA_izy & T==`Tfive & phi2)
			 | (OP==`ORA_zpx & T==`Tzero & phi1)
			 | (OP==`ORA_zpx & T==`Tzero & phi2)
			 | (OP==`ORA_zpx & T==`Tone & phi1)
			 | (OP==`ORA_zpx & T==`Tone & phi2)
			 | (OP==`ORA_zpx & T==`Ttwo & phi1)
			 | (OP==`ORA_zpx & T==`Ttwo & phi2)
			 | (OP==`ORA_zpx & T==`Tthree & phi1)
			 | (OP==`ORA_zpx & T==`Tthree & phi2)
			 | (OP==`ASL_zpx & T==`Tzero & phi1)
			 | (OP==`ASL_zpx & T==`Tzero & phi2)
			 | (OP==`ASL_zpx & T==`Tone & phi1)
			 | (OP==`ASL_zpx & T==`Tone & phi2)
			 | (OP==`ASL_zpx & T==`Ttwo & phi1)
			 | (OP==`ASL_zpx & T==`Ttwo & phi2)
			 | (OP==`ASL_zpx & T==`Tthree & phi1)
			 | (OP==`ASL_zpx & T==`Tthree & phi2)
			 | (OP==`ASL_zpx & T==`Tfour & phi1)
			 | (OP==`ASL_zpx & T==`Tfour & phi2)
			 | (OP==`ASL_zpx & T==`Tfive & phi1)
			 | (OP==`ASL_zpx & T==`Tfive & phi2)
			 | (OP==`CLC & T==`Tone & phi1)
			 | (OP==`CLC & T==`Tone & phi2)
			 | (OP==`CLC & T==`Ttwo & phi1)
			 | (OP==`CLC & T==`Ttwo & phi2)
			 | (OP==`ORA_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ORA_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`ORA_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`ORA_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`ORA_aby & T==`Tone & phi1)
			 | (OP==`ORA_aby & T==`Tone & phi2)
			 | (OP==`ORA_aby & T==`Ttwo & phi1)
			 | (OP==`ORA_aby & T==`Ttwo & phi2)
			 | (OP==`ORA_aby & T==`Tthree & phi1)
			 | (OP==`ORA_aby & T==`Tthree & phi2)
			 | (OP==`ORA_aby & T==`Tfour & phi1)
			 | (OP==`ORA_aby & T==`Tfour & phi2)
			 | (OP==`ORA_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ORA_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`ORA_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`ORA_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`ORA_abx & T==`Tone & phi1)
			 | (OP==`ORA_abx & T==`Tone & phi2)
			 | (OP==`ORA_abx & T==`Ttwo & phi1)
			 | (OP==`ORA_abx & T==`Ttwo & phi2)
			 | (OP==`ORA_abx & T==`Tthree & phi1)
			 | (OP==`ORA_abx & T==`Tthree & phi2)
			 | (OP==`ORA_abx & T==`Tfour & phi1)
			 | (OP==`ORA_abx & T==`Tfour & phi2)
			 | (OP==`ASL_abx & T==`Tzero & phi1)
			 | (OP==`ASL_abx & T==`Tzero & phi2)
			 | (OP==`ASL_abx & T==`Tone & phi1)
			 | (OP==`ASL_abx & T==`Tone & phi2)
			 | (OP==`ASL_abx & T==`Ttwo & phi1)
			 | (OP==`ASL_abx & T==`Ttwo & phi2)
			 | (OP==`ASL_abx & T==`Tthree & phi1)
			 | (OP==`ASL_abx & T==`Tthree & phi2)
			 | (OP==`ASL_abx & T==`Tfour & phi1)
			 | (OP==`ASL_abx & T==`Tfour & phi2)
			 | (OP==`ASL_abx & T==`Tfive & phi1)
			 | (OP==`ASL_abx & T==`Tfive & phi2)
			 | (OP==`ASL_abx & T==`Tsix & phi1)
			 | (OP==`ASL_abx & T==`Tsix & phi2)
			 | (OP==`JSR_abs & T==`Tzero & phi1)
			 | (OP==`JSR_abs & T==`Tzero & phi2)
			 | (OP==`JSR_abs & T==`Tone & phi1)
			 | (OP==`JSR_abs & T==`Tone & phi2)
			 | (OP==`JSR_abs & T==`Ttwo & phi1)
			 | (OP==`JSR_abs & T==`Ttwo & phi2)
			 | (OP==`JSR_abs & T==`Tthree & phi1)
			 | (OP==`JSR_abs & T==`Tthree & phi2)
			 | (OP==`JSR_abs & T==`Tfour & phi1)
			 | (OP==`JSR_abs & T==`Tfour & phi2)
			 | (OP==`JSR_abs & T==`Tfive & phi1)
			 | (OP==`JSR_abs & T==`Tfive & phi2)
			 | (OP==`AND_izx & T==`Tzero & phi1)
			 | (OP==`AND_izx & T==`Tzero & phi2)
			 | (OP==`AND_izx & T==`Tone & phi1)
			 | (OP==`AND_izx & T==`Tone & phi2)
			 | (OP==`AND_izx & T==`Ttwo & phi1)
			 | (OP==`AND_izx & T==`Ttwo & phi2)
			 | (OP==`AND_izx & T==`Tthree & phi1)
			 | (OP==`AND_izx & T==`Tthree & phi2)
			 | (OP==`AND_izx & T==`Tfour & phi1)
			 | (OP==`AND_izx & T==`Tfour & phi2)
			 | (OP==`AND_izx & T==`Tfive & phi1)
			 | (OP==`AND_izx & T==`Tfive & phi2)
			 | (OP==`BIT_zp & T==`Tzero & phi1)
			 | (OP==`BIT_zp & T==`Tzero & phi2)
			 | (OP==`BIT_zp & T==`Tone & phi1)
			 | (OP==`BIT_zp & T==`Tone & phi2)
			 | (OP==`BIT_zp & T==`Ttwo & phi1)
			 | (OP==`BIT_zp & T==`Ttwo & phi2)
			 | (OP==`AND_zp & T==`Tzero & phi1)
			 | (OP==`AND_zp & T==`Tzero & phi2)
			 | (OP==`AND_zp & T==`Tone & phi1)
			 | (OP==`AND_zp & T==`Tone & phi2)
			 | (OP==`AND_zp & T==`Ttwo & phi1)
			 | (OP==`AND_zp & T==`Ttwo & phi2)
			 | (OP==`ROL_zp & T==`Tzero & phi1)
			 | (OP==`ROL_zp & T==`Tzero & phi2)
			 | (OP==`ROL_zp & T==`Tone & phi1)
			 | (OP==`ROL_zp & T==`Tone & phi2)
			 | (OP==`ROL_zp & T==`Ttwo & phi1)
			 | (OP==`ROL_zp & T==`Ttwo & phi2)
			 | (OP==`ROL_zp & T==`Tthree & phi1)
			 | (OP==`ROL_zp & T==`Tthree & phi2)
			 | (OP==`ROL_zp & T==`Tfour & phi1)
			 | (OP==`ROL_zp & T==`Tfour & phi2)
			 | (OP==`PLP & T==`Tzero & phi1)
			 | (OP==`PLP & T==`Tzero & phi2)
			 | (OP==`PLP & T==`Tone & phi1)
			 | (OP==`PLP & T==`Tone & phi2)
			 | (OP==`PLP & T==`Ttwo & phi1)
			 | (OP==`PLP & T==`Ttwo & phi2)
			 | (OP==`PLP & T==`Tthree & phi1)
			 | (OP==`PLP & T==`Tthree & phi2)
			 | (OP==`AND_imm & T==`Tone & phi1)
			 | (OP==`AND_imm & T==`Tone & phi2)
			 | (OP==`AND_imm & T==`Ttwo & phi1)
			 | (OP==`AND_imm & T==`Ttwo & phi2)
			 | (OP==`ROL & T==`Tone & phi1)
			 | (OP==`ROL & T==`Tone & phi2)
			 | (OP==`ROL & T==`Ttwo & phi1)
			 | (OP==`ROL & T==`Ttwo & phi2)
			 | (OP==`BIT_abs & T==`Tzero & phi1)
			 | (OP==`BIT_abs & T==`Tzero & phi2)
			 | (OP==`BIT_abs & T==`Tone & phi1)
			 | (OP==`BIT_abs & T==`Tone & phi2)
			 | (OP==`BIT_abs & T==`Ttwo & phi1)
			 | (OP==`BIT_abs & T==`Ttwo & phi2)
			 | (OP==`BIT_abs & T==`Tthree & phi1)
			 | (OP==`BIT_abs & T==`Tthree & phi2)
			 | (OP==`AND_abs & T==`Tzero & phi1)
			 | (OP==`AND_abs & T==`Tzero & phi2)
			 | (OP==`AND_abs & T==`Tone & phi1)
			 | (OP==`AND_abs & T==`Tone & phi2)
			 | (OP==`AND_abs & T==`Ttwo & phi1)
			 | (OP==`AND_abs & T==`Ttwo & phi2)
			 | (OP==`AND_abs & T==`Tthree & phi1)
			 | (OP==`AND_abs & T==`Tthree & phi2)
			 | (OP==`ROL_abs & T==`Tzero & phi1)
			 | (OP==`ROL_abs & T==`Tzero & phi2)
			 | (OP==`ROL_abs & T==`Tone & phi1)
			 | (OP==`ROL_abs & T==`Tone & phi2)
			 | (OP==`ROL_abs & T==`Ttwo & phi1)
			 | (OP==`ROL_abs & T==`Ttwo & phi2)
			 | (OP==`ROL_abs & T==`Tthree & phi1)
			 | (OP==`ROL_abs & T==`Tthree & phi2)
			 | (OP==`ROL_abs & T==`Tfour & phi1)
			 | (OP==`ROL_abs & T==`Tfour & phi2)
			 | (OP==`ROL_abs & T==`Tfive & phi1)
			 | (OP==`ROL_abs & T==`Tfive & phi2)
			 | (OP==`BMI_rel & T==`Tzero & phi1)
			 | (OP==`BMI_rel & T==`Tzero & phi2)
			 | (OP==`BMI_rel & T==`Ttwo & phi1)
			 | (OP==`BMI_rel & T==`Ttwo & phi2)
			 | (OP==`BMI_rel & T==`Tthree & phi1)
			 | (OP==`BMI_rel & T==`Tthree & phi2)
			 | (OP==`BMI_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BMI_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BMI_rel & T==`T1BranchCross & phi1)
			 | (OP==`BMI_rel & T==`T1BranchCross & phi2)
			 | (OP==`BMI_rel & T==`T1NoBranch & phi1)
			 | (OP==`BMI_rel & T==`T1NoBranch & phi2)
			 | (OP==`AND_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`AND_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`AND_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`AND_izy & T==`TzeroCrossPg & phi2)
			 | (OP==`AND_izy & T==`Tone & phi1)
			 | (OP==`AND_izy & T==`Tone & phi2)
			 | (OP==`AND_izy & T==`Ttwo & phi1)
			 | (OP==`AND_izy & T==`Ttwo & phi2)
			 | (OP==`AND_izy & T==`Tthree & phi1)
			 | (OP==`AND_izy & T==`Tthree & phi2)
			 | (OP==`AND_izy & T==`Tfour & phi1)
			 | (OP==`AND_izy & T==`Tfour & phi2)
			 | (OP==`AND_izy & T==`Tfive & phi1)
			 | (OP==`AND_izy & T==`Tfive & phi2)
			 | (OP==`AND_zpx & T==`Tzero & phi1)
			 | (OP==`AND_zpx & T==`Tzero & phi2)
			 | (OP==`AND_zpx & T==`Tone & phi1)
			 | (OP==`AND_zpx & T==`Tone & phi2)
			 | (OP==`AND_zpx & T==`Ttwo & phi1)
			 | (OP==`AND_zpx & T==`Ttwo & phi2)
			 | (OP==`AND_zpx & T==`Tthree & phi1)
			 | (OP==`AND_zpx & T==`Tthree & phi2)
			 | (OP==`ROL_zpx & T==`Tzero & phi1)
			 | (OP==`ROL_zpx & T==`Tzero & phi2)
			 | (OP==`ROL_zpx & T==`Tone & phi1)
			 | (OP==`ROL_zpx & T==`Tone & phi2)
			 | (OP==`ROL_zpx & T==`Ttwo & phi1)
			 | (OP==`ROL_zpx & T==`Ttwo & phi2)
			 | (OP==`ROL_zpx & T==`Tthree & phi1)
			 | (OP==`ROL_zpx & T==`Tthree & phi2)
			 | (OP==`ROL_zpx & T==`Tfour & phi1)
			 | (OP==`ROL_zpx & T==`Tfour & phi2)
			 | (OP==`ROL_zpx & T==`Tfive & phi1)
			 | (OP==`ROL_zpx & T==`Tfive & phi2)
			 | (OP==`SEC & T==`Tone & phi1)
			 | (OP==`SEC & T==`Tone & phi2)
			 | (OP==`SEC & T==`Ttwo & phi1)
			 | (OP==`SEC & T==`Ttwo & phi2)
			 | (OP==`AND_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`AND_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`AND_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`AND_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`AND_aby & T==`Tone & phi1)
			 | (OP==`AND_aby & T==`Tone & phi2)
			 | (OP==`AND_aby & T==`Ttwo & phi1)
			 | (OP==`AND_aby & T==`Ttwo & phi2)
			 | (OP==`AND_aby & T==`Tthree & phi1)
			 | (OP==`AND_aby & T==`Tthree & phi2)
			 | (OP==`AND_aby & T==`Tfour & phi1)
			 | (OP==`AND_aby & T==`Tfour & phi2)
			 | (OP==`AND_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`AND_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`AND_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`AND_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`AND_abx & T==`Tone & phi1)
			 | (OP==`AND_abx & T==`Tone & phi2)
			 | (OP==`AND_abx & T==`Ttwo & phi1)
			 | (OP==`AND_abx & T==`Ttwo & phi2)
			 | (OP==`AND_abx & T==`Tthree & phi1)
			 | (OP==`AND_abx & T==`Tthree & phi2)
			 | (OP==`AND_abx & T==`Tfour & phi1)
			 | (OP==`AND_abx & T==`Tfour & phi2)
			 | (OP==`ROL_abx & T==`Tzero & phi1)
			 | (OP==`ROL_abx & T==`Tzero & phi2)
			 | (OP==`ROL_abx & T==`Tone & phi1)
			 | (OP==`ROL_abx & T==`Tone & phi2)
			 | (OP==`ROL_abx & T==`Ttwo & phi1)
			 | (OP==`ROL_abx & T==`Ttwo & phi2)
			 | (OP==`ROL_abx & T==`Tthree & phi1)
			 | (OP==`ROL_abx & T==`Tthree & phi2)
			 | (OP==`ROL_abx & T==`Tfour & phi1)
			 | (OP==`ROL_abx & T==`Tfour & phi2)
			 | (OP==`ROL_abx & T==`Tfive & phi1)
			 | (OP==`ROL_abx & T==`Tfive & phi2)
			 | (OP==`ROL_abx & T==`Tsix & phi1)
			 | (OP==`ROL_abx & T==`Tsix & phi2)
			 | (OP==`RTI & T==`Tzero & phi1)
			 | (OP==`RTI & T==`Tzero & phi2)
			 | (OP==`RTI & T==`Tone & phi1)
			 | (OP==`RTI & T==`Tone & phi2)
			 | (OP==`RTI & T==`Ttwo & phi1)
			 | (OP==`RTI & T==`Ttwo & phi2)
			 | (OP==`RTI & T==`Tthree & phi1)
			 | (OP==`RTI & T==`Tthree & phi2)
			 | (OP==`RTI & T==`Tfour & phi1)
			 | (OP==`RTI & T==`Tfour & phi2)
			 | (OP==`RTI & T==`Tfive & phi1)
			 | (OP==`RTI & T==`Tfive & phi2)
			 | (OP==`EOR_izx & T==`Tzero & phi1)
			 | (OP==`EOR_izx & T==`Tzero & phi2)
			 | (OP==`EOR_izx & T==`Tone & phi1)
			 | (OP==`EOR_izx & T==`Tone & phi2)
			 | (OP==`EOR_izx & T==`Ttwo & phi1)
			 | (OP==`EOR_izx & T==`Ttwo & phi2)
			 | (OP==`EOR_izx & T==`Tthree & phi1)
			 | (OP==`EOR_izx & T==`Tthree & phi2)
			 | (OP==`EOR_izx & T==`Tfour & phi1)
			 | (OP==`EOR_izx & T==`Tfour & phi2)
			 | (OP==`EOR_izx & T==`Tfive & phi1)
			 | (OP==`EOR_izx & T==`Tfive & phi2)
			 | (OP==`EOR_zp & T==`Tzero & phi1)
			 | (OP==`EOR_zp & T==`Tzero & phi2)
			 | (OP==`EOR_zp & T==`Tone & phi1)
			 | (OP==`EOR_zp & T==`Tone & phi2)
			 | (OP==`EOR_zp & T==`Ttwo & phi1)
			 | (OP==`EOR_zp & T==`Ttwo & phi2)
			 | (OP==`LSR_zp & T==`Tzero & phi1)
			 | (OP==`LSR_zp & T==`Tzero & phi2)
			 | (OP==`LSR_zp & T==`Tone & phi1)
			 | (OP==`LSR_zp & T==`Tone & phi2)
			 | (OP==`LSR_zp & T==`Ttwo & phi1)
			 | (OP==`LSR_zp & T==`Ttwo & phi2)
			 | (OP==`LSR_zp & T==`Tthree & phi1)
			 | (OP==`LSR_zp & T==`Tthree & phi2)
			 | (OP==`LSR_zp & T==`Tfour & phi1)
			 | (OP==`LSR_zp & T==`Tfour & phi2)
			 | (OP==`PHA & T==`Tzero & phi1)
			 | (OP==`PHA & T==`Tzero & phi2)
			 | (OP==`PHA & T==`Tone & phi1)
			 | (OP==`PHA & T==`Tone & phi2)
			 | (OP==`PHA & T==`Ttwo & phi1)
			 | (OP==`PHA & T==`Ttwo & phi2)
			 | (OP==`EOR_imm & T==`Tone & phi1)
			 | (OP==`EOR_imm & T==`Tone & phi2)
			 | (OP==`EOR_imm & T==`Ttwo & phi1)
			 | (OP==`EOR_imm & T==`Ttwo & phi2)
			 | (OP==`LSR & T==`Tone & phi1)
			 | (OP==`LSR & T==`Tone & phi2)
			 | (OP==`LSR & T==`Ttwo & phi1)
			 | (OP==`LSR & T==`Ttwo & phi2)
			 | (OP==`JMP_abs & T==`Tzero & phi1)
			 | (OP==`JMP_abs & T==`Tzero & phi2)
			 | (OP==`JMP_abs & T==`Tone & phi1)
			 | (OP==`JMP_abs & T==`Tone & phi2)
			 | (OP==`JMP_abs & T==`Ttwo & phi1)
			 | (OP==`JMP_abs & T==`Ttwo & phi2)
			 | (OP==`EOR_abs & T==`Tzero & phi1)
			 | (OP==`EOR_abs & T==`Tzero & phi2)
			 | (OP==`EOR_abs & T==`Tone & phi1)
			 | (OP==`EOR_abs & T==`Tone & phi2)
			 | (OP==`EOR_abs & T==`Ttwo & phi1)
			 | (OP==`EOR_abs & T==`Ttwo & phi2)
			 | (OP==`EOR_abs & T==`Tthree & phi1)
			 | (OP==`EOR_abs & T==`Tthree & phi2)
			 | (OP==`LSR_abs & T==`Tzero & phi1)
			 | (OP==`LSR_abs & T==`Tzero & phi2)
			 | (OP==`LSR_abs & T==`Tone & phi1)
			 | (OP==`LSR_abs & T==`Tone & phi2)
			 | (OP==`LSR_abs & T==`Ttwo & phi1)
			 | (OP==`LSR_abs & T==`Ttwo & phi2)
			 | (OP==`LSR_abs & T==`Tthree & phi1)
			 | (OP==`LSR_abs & T==`Tthree & phi2)
			 | (OP==`LSR_abs & T==`Tfour & phi1)
			 | (OP==`LSR_abs & T==`Tfour & phi2)
			 | (OP==`LSR_abs & T==`Tfive & phi1)
			 | (OP==`LSR_abs & T==`Tfive & phi2)
			 | (OP==`BVC_rel & T==`Tzero & phi1)
			 | (OP==`BVC_rel & T==`Tzero & phi2)
			 | (OP==`BVC_rel & T==`Ttwo & phi1)
			 | (OP==`BVC_rel & T==`Ttwo & phi2)
			 | (OP==`BVC_rel & T==`Tthree & phi1)
			 | (OP==`BVC_rel & T==`Tthree & phi2)
			 | (OP==`BVC_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BVC_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BVC_rel & T==`T1BranchCross & phi1)
			 | (OP==`BVC_rel & T==`T1BranchCross & phi2)
			 | (OP==`BVC_rel & T==`T1NoBranch & phi1)
			 | (OP==`BVC_rel & T==`T1NoBranch & phi2)
			 | (OP==`EOR_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`EOR_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`EOR_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`EOR_izy & T==`TzeroCrossPg & phi2)
			 | (OP==`EOR_izy & T==`Tone & phi1)
			 | (OP==`EOR_izy & T==`Tone & phi2)
			 | (OP==`EOR_izy & T==`Ttwo & phi1)
			 | (OP==`EOR_izy & T==`Ttwo & phi2)
			 | (OP==`EOR_izy & T==`Tthree & phi1)
			 | (OP==`EOR_izy & T==`Tthree & phi2)
			 | (OP==`EOR_izy & T==`Tfour & phi1)
			 | (OP==`EOR_izy & T==`Tfour & phi2)
			 | (OP==`EOR_izy & T==`Tfive & phi1)
			 | (OP==`EOR_izy & T==`Tfive & phi2)
			 | (OP==`EOR_zpx & T==`Tzero & phi1)
			 | (OP==`EOR_zpx & T==`Tzero & phi2)
			 | (OP==`EOR_zpx & T==`Tone & phi1)
			 | (OP==`EOR_zpx & T==`Tone & phi2)
			 | (OP==`EOR_zpx & T==`Ttwo & phi1)
			 | (OP==`EOR_zpx & T==`Ttwo & phi2)
			 | (OP==`EOR_zpx & T==`Tthree & phi1)
			 | (OP==`EOR_zpx & T==`Tthree & phi2)
			 | (OP==`LSR_zpx & T==`Tzero & phi1)
			 | (OP==`LSR_zpx & T==`Tzero & phi2)
			 | (OP==`LSR_zpx & T==`Tone & phi1)
			 | (OP==`LSR_zpx & T==`Tone & phi2)
			 | (OP==`LSR_zpx & T==`Ttwo & phi1)
			 | (OP==`LSR_zpx & T==`Ttwo & phi2)
			 | (OP==`LSR_zpx & T==`Tthree & phi1)
			 | (OP==`LSR_zpx & T==`Tthree & phi2)
			 | (OP==`LSR_zpx & T==`Tfour & phi1)
			 | (OP==`LSR_zpx & T==`Tfour & phi2)
			 | (OP==`LSR_zpx & T==`Tfive & phi1)
			 | (OP==`LSR_zpx & T==`Tfive & phi2)
			 | (OP==`CLI & T==`Tone & phi1)
			 | (OP==`CLI & T==`Tone & phi2)
			 | (OP==`CLI & T==`Ttwo & phi1)
			 | (OP==`CLI & T==`Ttwo & phi2)
			 | (OP==`EOR_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`EOR_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`EOR_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`EOR_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`EOR_aby & T==`Tone & phi1)
			 | (OP==`EOR_aby & T==`Tone & phi2)
			 | (OP==`EOR_aby & T==`Ttwo & phi1)
			 | (OP==`EOR_aby & T==`Ttwo & phi2)
			 | (OP==`EOR_aby & T==`Tthree & phi1)
			 | (OP==`EOR_aby & T==`Tthree & phi2)
			 | (OP==`EOR_aby & T==`Tfour & phi1)
			 | (OP==`EOR_aby & T==`Tfour & phi2)
			 | (OP==`EOR_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`EOR_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`EOR_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`EOR_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`EOR_abx & T==`Tone & phi1)
			 | (OP==`EOR_abx & T==`Tone & phi2)
			 | (OP==`EOR_abx & T==`Ttwo & phi1)
			 | (OP==`EOR_abx & T==`Ttwo & phi2)
			 | (OP==`EOR_abx & T==`Tthree & phi1)
			 | (OP==`EOR_abx & T==`Tthree & phi2)
			 | (OP==`EOR_abx & T==`Tfour & phi1)
			 | (OP==`EOR_abx & T==`Tfour & phi2)
			 | (OP==`LSR_abx & T==`Tzero & phi1)
			 | (OP==`LSR_abx & T==`Tzero & phi2)
			 | (OP==`LSR_abx & T==`Tone & phi1)
			 | (OP==`LSR_abx & T==`Tone & phi2)
			 | (OP==`LSR_abx & T==`Ttwo & phi1)
			 | (OP==`LSR_abx & T==`Ttwo & phi2)
			 | (OP==`LSR_abx & T==`Tthree & phi1)
			 | (OP==`LSR_abx & T==`Tthree & phi2)
			 | (OP==`LSR_abx & T==`Tfour & phi1)
			 | (OP==`LSR_abx & T==`Tfour & phi2)
			 | (OP==`LSR_abx & T==`Tfive & phi1)
			 | (OP==`LSR_abx & T==`Tfive & phi2)
			 | (OP==`LSR_abx & T==`Tsix & phi1)
			 | (OP==`LSR_abx & T==`Tsix & phi2)
			 | (OP==`RTS & T==`Tzero & phi1)
			 | (OP==`RTS & T==`Tzero & phi2)
			 | (OP==`RTS & T==`Tone & phi1)
			 | (OP==`RTS & T==`Tone & phi2)
			 | (OP==`RTS & T==`Ttwo & phi1)
			 | (OP==`RTS & T==`Ttwo & phi2)
			 | (OP==`RTS & T==`Tthree & phi1)
			 | (OP==`RTS & T==`Tthree & phi2)
			 | (OP==`RTS & T==`Tfour & phi1)
			 | (OP==`RTS & T==`Tfour & phi2)
			 | (OP==`RTS & T==`Tfive & phi1)
			 | (OP==`RTS & T==`Tfive & phi2)
			 | (OP==`ADC_izx & T==`Tzero & phi1)
			 | (OP==`ADC_izx & T==`Tzero & phi2)
			 | (OP==`ADC_izx & T==`Tone & phi1 & !decMode)
			 | (OP==`ADC_izx & T==`Tone & phi2 & !decMode)
			 | (OP==`ADC_izx & T==`Ttwo & phi1)
			 | (OP==`ADC_izx & T==`Ttwo & phi2)
			 | (OP==`ADC_izx & T==`Tthree & phi1)
			 | (OP==`ADC_izx & T==`Tthree & phi2)
			 | (OP==`ADC_izx & T==`Tfour & phi1)
			 | (OP==`ADC_izx & T==`Tfour & phi2)
			 | (OP==`ADC_izx & T==`Tfive & phi1)
			 | (OP==`ADC_izx & T==`Tfive & phi2)
			 | (OP==`ADC_zp & T==`Tzero & phi1)
			 | (OP==`ADC_zp & T==`Tzero & phi2)
			 | (OP==`ADC_zp & T==`Tone & phi1 & !decMode)
			 | (OP==`ADC_zp & T==`Tone & phi2 & !decMode)
			 | (OP==`ADC_zp & T==`Ttwo & phi1)
			 | (OP==`ADC_zp & T==`Ttwo & phi2)
			 | (OP==`ROR_zp & T==`Tzero & phi1)
			 | (OP==`ROR_zp & T==`Tzero & phi2)
			 | (OP==`ROR_zp & T==`Tone & phi1)
			 | (OP==`ROR_zp & T==`Tone & phi2)
			 | (OP==`ROR_zp & T==`Ttwo & phi1)
			 | (OP==`ROR_zp & T==`Ttwo & phi2)
			 | (OP==`ROR_zp & T==`Tthree & phi1)
			 | (OP==`ROR_zp & T==`Tthree & phi2)
			 | (OP==`ROR_zp & T==`Tfour & phi1)
			 | (OP==`ROR_zp & T==`Tfour & phi2)
			 | (OP==`PLA & T==`Tzero & phi1)
			 | (OP==`PLA & T==`Tzero & phi2)
			 | (OP==`PLA & T==`Tone & phi1)
			 | (OP==`PLA & T==`Tone & phi2)
			 | (OP==`PLA & T==`Ttwo & phi1)
			 | (OP==`PLA & T==`Ttwo & phi2)
			 | (OP==`PLA & T==`Tthree & phi1)
			 | (OP==`PLA & T==`Tthree & phi2)
			 | (OP==`ADC_imm & T==`Tone & phi1 & !decMode)
			 | (OP==`ADC_imm & T==`Tone & phi2 & !decMode)
			 | (OP==`ADC_imm & T==`Ttwo & phi1)
			 | (OP==`ADC_imm & T==`Ttwo & phi2)
			 | (OP==`ROR & T==`Tone & phi1)
			 | (OP==`ROR & T==`Tone & phi2)
			 | (OP==`ROR & T==`Ttwo & phi1)
			 | (OP==`ROR & T==`Ttwo & phi2)
			 | (OP==`JMP_zp & T==`Tzero & phi1)
			 | (OP==`JMP_zp & T==`Tzero & phi2)
			 | (OP==`JMP_zp & T==`Tone & phi1)
			 | (OP==`JMP_zp & T==`Tone & phi2)
			 | (OP==`JMP_zp & T==`Ttwo & phi1)
			 | (OP==`JMP_zp & T==`Ttwo & phi2)
			 | (OP==`JMP_zp & T==`Tthree & phi1)
			 | (OP==`JMP_zp & T==`Tthree & phi2)
			 | (OP==`JMP_zp & T==`Tfour & phi1)
			 | (OP==`JMP_zp & T==`Tfour & phi2)
			 | (OP==`ADC_abs & T==`Tzero & phi1)
			 | (OP==`ADC_abs & T==`Tzero & phi2)
			 | (OP==`ADC_abs & T==`Tone & phi1 & !decMode)
			 | (OP==`ADC_abs & T==`Tone & phi2 & !decMode)
			 | (OP==`ADC_abs & T==`Ttwo & phi1)
			 | (OP==`ADC_abs & T==`Ttwo & phi2)
			 | (OP==`ADC_abs & T==`Tthree & phi1)
			 | (OP==`ADC_abs & T==`Tthree & phi2)
			 | (OP==`ROR_abs & T==`Tzero & phi1)
			 | (OP==`ROR_abs & T==`Tzero & phi2)
			 | (OP==`ROR_abs & T==`Tone & phi1)
			 | (OP==`ROR_abs & T==`Tone & phi2)
			 | (OP==`ROR_abs & T==`Ttwo & phi1)
			 | (OP==`ROR_abs & T==`Ttwo & phi2)
			 | (OP==`ROR_abs & T==`Tthree & phi1)
			 | (OP==`ROR_abs & T==`Tthree & phi2)
			 | (OP==`ROR_abs & T==`Tfour & phi1)
			 | (OP==`ROR_abs & T==`Tfour & phi2)
			 | (OP==`ROR_abs & T==`Tfive & phi1)
			 | (OP==`ROR_abs & T==`Tfive & phi2)
			 | (OP==`BVS_rel & T==`Tzero & phi1)
			 | (OP==`BVS_rel & T==`Tzero & phi2)
			 | (OP==`BVS_rel & T==`Ttwo & phi1)
			 | (OP==`BVS_rel & T==`Ttwo & phi2)
			 | (OP==`BVS_rel & T==`Tthree & phi1)
			 | (OP==`BVS_rel & T==`Tthree & phi2)
			 | (OP==`BVS_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BVS_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BVS_rel & T==`T1BranchCross & phi1)
			 | (OP==`BVS_rel & T==`T1BranchCross & phi2)
			 | (OP==`BVS_rel & T==`T1NoBranch & phi1)
			 | (OP==`BVS_rel & T==`T1NoBranch & phi2)
			 | (OP==`ADC_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ADC_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`ADC_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`ADC_izy & T==`TzeroCrossPg & phi2)
			 | (OP==`ADC_izy & T==`Tone & phi1 & !decMode)
			 | (OP==`ADC_izy & T==`Tone & phi2 & !decMode)
			 | (OP==`ADC_izy & T==`Ttwo & phi1)
			 | (OP==`ADC_izy & T==`Ttwo & phi2)
			 | (OP==`ADC_izy & T==`Tthree & phi1)
			 | (OP==`ADC_izy & T==`Tthree & phi2)
			 | (OP==`ADC_izy & T==`Tfour & phi1)
			 | (OP==`ADC_izy & T==`Tfour & phi2)
			 | (OP==`ADC_izy & T==`Tfive & phi1)
			 | (OP==`ADC_izy & T==`Tfive & phi2)
			 | (OP==`ADC_zpx & T==`Tzero & phi1)
			 | (OP==`ADC_zpx & T==`Tzero & phi2)
			 | (OP==`ADC_zpx & T==`Tone & phi1 & !decMode)
			 | (OP==`ADC_zpx & T==`Tone & phi2 & !decMode)
			 | (OP==`ADC_zpx & T==`Ttwo & phi1)
			 | (OP==`ADC_zpx & T==`Ttwo & phi2)
			 | (OP==`ADC_zpx & T==`Tthree & phi1)
			 | (OP==`ADC_zpx & T==`Tthree & phi2)
			 | (OP==`ROR_zpx & T==`Tzero & phi1)
			 | (OP==`ROR_zpx & T==`Tzero & phi2)
			 | (OP==`ROR_zpx & T==`Tone & phi1)
			 | (OP==`ROR_zpx & T==`Tone & phi2)
			 | (OP==`ROR_zpx & T==`Ttwo & phi1)
			 | (OP==`ROR_zpx & T==`Ttwo & phi2)
			 | (OP==`ROR_zpx & T==`Tthree & phi1)
			 | (OP==`ROR_zpx & T==`Tthree & phi2)
			 | (OP==`ROR_zpx & T==`Tfour & phi1)
			 | (OP==`ROR_zpx & T==`Tfour & phi2)
			 | (OP==`ROR_zpx & T==`Tfive & phi1)
			 | (OP==`ROR_zpx & T==`Tfive & phi2)
			 | (OP==`SEI & T==`Tone & phi1)
			 | (OP==`SEI & T==`Tone & phi2)
			 | (OP==`SEI & T==`Ttwo & phi1)
			 | (OP==`SEI & T==`Ttwo & phi2)
			 | (OP==`ADC_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ADC_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`ADC_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`ADC_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`ADC_aby & T==`Tone & phi1 & !decMode)
			 | (OP==`ADC_aby & T==`Tone & phi2 & !decMode)
			 | (OP==`ADC_aby & T==`Ttwo & phi1)
			 | (OP==`ADC_aby & T==`Ttwo & phi2)
			 | (OP==`ADC_aby & T==`Tthree & phi1)
			 | (OP==`ADC_aby & T==`Tthree & phi2)
			 | (OP==`ADC_aby & T==`Tfour & phi1)
			 | (OP==`ADC_aby & T==`Tfour & phi2)
			 | (OP==`ADC_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ADC_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`ADC_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`ADC_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`ADC_abx & T==`Tone & phi1 & !decMode)
			 | (OP==`ADC_abx & T==`Tone & phi2 & !decMode)
			 | (OP==`ADC_abx & T==`Ttwo & phi1)
			 | (OP==`ADC_abx & T==`Ttwo & phi2)
			 | (OP==`ADC_abx & T==`Tthree & phi1)
			 | (OP==`ADC_abx & T==`Tthree & phi2)
			 | (OP==`ADC_abx & T==`Tfour & phi1)
			 | (OP==`ADC_abx & T==`Tfour & phi2)
			 | (OP==`ROR_abx & T==`Tzero & phi1)
			 | (OP==`ROR_abx & T==`Tzero & phi2)
			 | (OP==`ROR_abx & T==`Tone & phi1)
			 | (OP==`ROR_abx & T==`Tone & phi2)
			 | (OP==`ROR_abx & T==`Ttwo & phi1)
			 | (OP==`ROR_abx & T==`Ttwo & phi2)
			 | (OP==`ROR_abx & T==`Tthree & phi1)
			 | (OP==`ROR_abx & T==`Tthree & phi2)
			 | (OP==`ROR_abx & T==`Tfour & phi1)
			 | (OP==`ROR_abx & T==`Tfour & phi2)
			 | (OP==`ROR_abx & T==`Tfive & phi1)
			 | (OP==`ROR_abx & T==`Tfive & phi2)
			 | (OP==`ROR_abx & T==`Tsix & phi1)
			 | (OP==`ROR_abx & T==`Tsix & phi2)
			 | (OP==`STA_izx & T==`Tzero & phi1)
			 | (OP==`STA_izx & T==`Tzero & phi2)
			 | (OP==`STA_izx & T==`Tone & phi1)
			 | (OP==`STA_izx & T==`Tone & phi2)
			 | (OP==`STA_izx & T==`Ttwo & phi1)
			 | (OP==`STA_izx & T==`Ttwo & phi2)
			 | (OP==`STA_izx & T==`Tthree & phi1)
			 | (OP==`STA_izx & T==`Tthree & phi2)
			 | (OP==`STA_izx & T==`Tfour & phi1)
			 | (OP==`STA_izx & T==`Tfour & phi2)
			 | (OP==`STA_izx & T==`Tfive & phi1)
			 | (OP==`STA_izx & T==`Tfive & phi2)
			 | (OP==`STY_zp & T==`Tzero & phi1)
			 | (OP==`STY_zp & T==`Tzero & phi2)
			 | (OP==`STY_zp & T==`Tone & phi1)
			 | (OP==`STY_zp & T==`Tone & phi2)
			 | (OP==`STY_zp & T==`Ttwo & phi1)
			 | (OP==`STY_zp & T==`Ttwo & phi2)
			 | (OP==`STA_zp & T==`Tzero & phi1)
			 | (OP==`STA_zp & T==`Tzero & phi2)
			 | (OP==`STA_zp & T==`Tone & phi1)
			 | (OP==`STA_zp & T==`Tone & phi2)
			 | (OP==`STA_zp & T==`Ttwo & phi1)
			 | (OP==`STA_zp & T==`Ttwo & phi2)
			 | (OP==`STX_zp & T==`Tzero & phi1)
			 | (OP==`STX_zp & T==`Tzero & phi2)
			 | (OP==`STX_zp & T==`Tone & phi1)
			 | (OP==`STX_zp & T==`Tone & phi2)
			 | (OP==`STX_zp & T==`Ttwo & phi1)
			 | (OP==`STX_zp & T==`Ttwo & phi2)
			 | (OP==`DEY & T==`Tone & phi1)
			 | (OP==`DEY & T==`Tone & phi2)
			 | (OP==`DEY & T==`Ttwo & phi1)
			 | (OP==`DEY & T==`Ttwo & phi2)
			 | (OP==`TXA & T==`Tone & phi1)
			 | (OP==`TXA & T==`Tone & phi2)
			 | (OP==`TXA & T==`Ttwo & phi1)
			 | (OP==`TXA & T==`Ttwo & phi2)
			 | (OP==`STY_abs & T==`Tzero & phi1)
			 | (OP==`STY_abs & T==`Tzero & phi2)
			 | (OP==`STY_abs & T==`Tone & phi1)
			 | (OP==`STY_abs & T==`Tone & phi2)
			 | (OP==`STY_abs & T==`Ttwo & phi1)
			 | (OP==`STY_abs & T==`Ttwo & phi2)
			 | (OP==`STY_abs & T==`Tthree & phi1)
			 | (OP==`STY_abs & T==`Tthree & phi2)
			 | (OP==`STA_abs & T==`Tzero & phi1)
			 | (OP==`STA_abs & T==`Tzero & phi2)
			 | (OP==`STA_abs & T==`Tone & phi1)
			 | (OP==`STA_abs & T==`Tone & phi2)
			 | (OP==`STA_abs & T==`Ttwo & phi1)
			 | (OP==`STA_abs & T==`Ttwo & phi2)
			 | (OP==`STA_abs & T==`Tthree & phi1)
			 | (OP==`STA_abs & T==`Tthree & phi2)
			 | (OP==`STX_abs & T==`Tzero & phi1)
			 | (OP==`STX_abs & T==`Tzero & phi2)
			 | (OP==`STX_abs & T==`Tone & phi1)
			 | (OP==`STX_abs & T==`Tone & phi2)
			 | (OP==`STX_abs & T==`Ttwo & phi1)
			 | (OP==`STX_abs & T==`Ttwo & phi2)
			 | (OP==`STX_abs & T==`Tthree & phi1)
			 | (OP==`STX_abs & T==`Tthree & phi2)
			 | (OP==`BCC_rel & T==`Tzero & phi1)
			 | (OP==`BCC_rel & T==`Tzero & phi2)
			 | (OP==`BCC_rel & T==`Ttwo & phi1)
			 | (OP==`BCC_rel & T==`Ttwo & phi2)
			 | (OP==`BCC_rel & T==`Tthree & phi1)
			 | (OP==`BCC_rel & T==`Tthree & phi2)
			 | (OP==`BCC_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BCC_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BCC_rel & T==`T1BranchCross & phi1)
			 | (OP==`BCC_rel & T==`T1BranchCross & phi2)
			 | (OP==`BCC_rel & T==`T1NoBranch & phi1)
			 | (OP==`BCC_rel & T==`T1NoBranch & phi2)
			 | (OP==`STA_izy & T==`Tzero & phi1)
			 | (OP==`STA_izy & T==`Tzero & phi2)
			 | (OP==`STA_izy & T==`Tone & phi1)
			 | (OP==`STA_izy & T==`Tone & phi2)
			 | (OP==`STA_izy & T==`Ttwo & phi1)
			 | (OP==`STA_izy & T==`Ttwo & phi2)
			 | (OP==`STA_izy & T==`Tthree & phi1)
			 | (OP==`STA_izy & T==`Tthree & phi2)
			 | (OP==`STA_izy & T==`Tfour & phi1)
			 | (OP==`STA_izy & T==`Tfour & phi2)
			 | (OP==`STA_izy & T==`Tfive & phi1)
			 | (OP==`STA_izy & T==`Tfive & phi2)
			 | (OP==`STY_zpx & T==`Tzero & phi1)
			 | (OP==`STY_zpx & T==`Tzero & phi2)
			 | (OP==`STY_zpx & T==`Tone & phi1)
			 | (OP==`STY_zpx & T==`Tone & phi2)
			 | (OP==`STY_zpx & T==`Ttwo & phi1)
			 | (OP==`STY_zpx & T==`Ttwo & phi2)
			 | (OP==`STY_zpx & T==`Tthree & phi1)
			 | (OP==`STY_zpx & T==`Tthree & phi2)
			 | (OP==`STA_zpx & T==`Tzero & phi1)
			 | (OP==`STA_zpx & T==`Tzero & phi2)
			 | (OP==`STA_zpx & T==`Tone & phi1)
			 | (OP==`STA_zpx & T==`Tone & phi2)
			 | (OP==`STA_zpx & T==`Ttwo & phi1)
			 | (OP==`STA_zpx & T==`Ttwo & phi2)
			 | (OP==`STA_zpx & T==`Tthree & phi1)
			 | (OP==`STA_zpx & T==`Tthree & phi2)
			 | (OP==`STX_zpy & T==`Tzero & phi1)
			 | (OP==`STX_zpy & T==`Tzero & phi2)
			 | (OP==`STX_zpy & T==`Tone & phi1)
			 | (OP==`STX_zpy & T==`Tone & phi2)
			 | (OP==`STX_zpy & T==`Ttwo & phi1)
			 | (OP==`STX_zpy & T==`Ttwo & phi2)
			 | (OP==`STX_zpy & T==`Tthree & phi1)
			 | (OP==`STX_zpy & T==`Tthree & phi2)
			 | (OP==`TYA & T==`Tone & phi1)
			 | (OP==`TYA & T==`Tone & phi2)
			 | (OP==`TYA & T==`Ttwo & phi1)
			 | (OP==`TYA & T==`Ttwo & phi2)
			 | (OP==`STA_aby & T==`Tzero & phi1)
			 | (OP==`STA_aby & T==`Tzero & phi2)
			 | (OP==`STA_aby & T==`Tone & phi1)
			 | (OP==`STA_aby & T==`Tone & phi2)
			 | (OP==`STA_aby & T==`Ttwo & phi1)
			 | (OP==`STA_aby & T==`Ttwo & phi2)
			 | (OP==`STA_aby & T==`Tthree & phi1)
			 | (OP==`STA_aby & T==`Tthree & phi2)
			 | (OP==`STA_aby & T==`Tfour & phi1)
			 | (OP==`STA_aby & T==`Tfour & phi2)
			 | (OP==`TXS & T==`Tone & phi1)
			 | (OP==`TXS & T==`Tone & phi2)
			 | (OP==`TXS & T==`Ttwo & phi1)
			 | (OP==`TXS & T==`Ttwo & phi2)
			 | (OP==`STA_abx & T==`Tzero & phi1)
			 | (OP==`STA_abx & T==`Tzero & phi2)
			 | (OP==`STA_abx & T==`Tone & phi1)
			 | (OP==`STA_abx & T==`Tone & phi2)
			 | (OP==`STA_abx & T==`Ttwo & phi1)
			 | (OP==`STA_abx & T==`Ttwo & phi2)
			 | (OP==`STA_abx & T==`Tthree & phi1)
			 | (OP==`STA_abx & T==`Tthree & phi2)
			 | (OP==`STA_abx & T==`Tfour & phi1)
			 | (OP==`STA_abx & T==`Tfour & phi2)
			 | (OP==`LDY_imm & T==`Tone & phi1)
			 | (OP==`LDY_imm & T==`Tone & phi2)
			 | (OP==`LDY_imm & T==`Ttwo & phi1)
			 | (OP==`LDY_imm & T==`Ttwo & phi2)
			 | (OP==`LDA_izx & T==`Tzero & phi1)
			 | (OP==`LDA_izx & T==`Tzero & phi2)
			 | (OP==`LDA_izx & T==`Tone & phi1)
			 | (OP==`LDA_izx & T==`Tone & phi2)
			 | (OP==`LDA_izx & T==`Ttwo & phi1)
			 | (OP==`LDA_izx & T==`Ttwo & phi2)
			 | (OP==`LDA_izx & T==`Tthree & phi1)
			 | (OP==`LDA_izx & T==`Tthree & phi2)
			 | (OP==`LDA_izx & T==`Tfour & phi1)
			 | (OP==`LDA_izx & T==`Tfour & phi2)
			 | (OP==`LDA_izx & T==`Tfive & phi1)
			 | (OP==`LDA_izx & T==`Tfive & phi2)
			 | (OP==`LDX_imm & T==`Tone & phi1)
			 | (OP==`LDX_imm & T==`Tone & phi2)
			 | (OP==`LDX_imm & T==`Ttwo & phi1)
			 | (OP==`LDX_imm & T==`Ttwo & phi2)
			 | (OP==`LDY_zp & T==`Tzero & phi1)
			 | (OP==`LDY_zp & T==`Tzero & phi2)
			 | (OP==`LDY_zp & T==`Tone & phi1)
			 | (OP==`LDY_zp & T==`Tone & phi2)
			 | (OP==`LDY_zp & T==`Ttwo & phi1)
			 | (OP==`LDY_zp & T==`Ttwo & phi2)
			 | (OP==`LDA_zp & T==`Tzero & phi1)
			 | (OP==`LDA_zp & T==`Tzero & phi2)
			 | (OP==`LDA_zp & T==`Tone & phi1)
			 | (OP==`LDA_zp & T==`Tone & phi2)
			 | (OP==`LDA_zp & T==`Ttwo & phi1)
			 | (OP==`LDA_zp & T==`Ttwo & phi2)
			 | (OP==`LDX_zp & T==`Tzero & phi1)
			 | (OP==`LDX_zp & T==`Tzero & phi2)
			 | (OP==`LDX_zp & T==`Tone & phi1)
			 | (OP==`LDX_zp & T==`Tone & phi2)
			 | (OP==`LDX_zp & T==`Ttwo & phi1)
			 | (OP==`LDX_zp & T==`Ttwo & phi2)
			 | (OP==`TAY & T==`Tone & phi1)
			 | (OP==`TAY & T==`Tone & phi2)
			 | (OP==`TAY & T==`Ttwo & phi1)
			 | (OP==`TAY & T==`Ttwo & phi2)
			 | (OP==`LDA_imm & T==`Tone & phi1)
			 | (OP==`LDA_imm & T==`Tone & phi2)
			 | (OP==`LDA_imm & T==`Ttwo & phi1)
			 | (OP==`LDA_imm & T==`Ttwo & phi2)
			 | (OP==`TAX & T==`Tone & phi1)
			 | (OP==`TAX & T==`Tone & phi2)
			 | (OP==`TAX & T==`Ttwo & phi1)
			 | (OP==`TAX & T==`Ttwo & phi2)
			 | (OP==`LDY_abs & T==`Tzero & phi1)
			 | (OP==`LDY_abs & T==`Tzero & phi2)
			 | (OP==`LDY_abs & T==`Tone & phi1)
			 | (OP==`LDY_abs & T==`Tone & phi2)
			 | (OP==`LDY_abs & T==`Ttwo & phi1)
			 | (OP==`LDY_abs & T==`Ttwo & phi2)
			 | (OP==`LDY_abs & T==`Tthree & phi1)
			 | (OP==`LDY_abs & T==`Tthree & phi2)
			 | (OP==`LDA_abs & T==`Tzero & phi1)
			 | (OP==`LDA_abs & T==`Tzero & phi2)
			 | (OP==`LDA_abs & T==`Tone & phi1)
			 | (OP==`LDA_abs & T==`Tone & phi2)
			 | (OP==`LDA_abs & T==`Ttwo & phi1)
			 | (OP==`LDA_abs & T==`Ttwo & phi2)
			 | (OP==`LDA_abs & T==`Tthree & phi1)
			 | (OP==`LDA_abs & T==`Tthree & phi2)
			 | (OP==`LDX_abs & T==`Tzero & phi1)
			 | (OP==`LDX_abs & T==`Tzero & phi2)
			 | (OP==`LDX_abs & T==`Tone & phi1)
			 | (OP==`LDX_abs & T==`Tone & phi2)
			 | (OP==`LDX_abs & T==`Ttwo & phi1)
			 | (OP==`LDX_abs & T==`Ttwo & phi2)
			 | (OP==`LDX_abs & T==`Tthree & phi1)
			 | (OP==`LDX_abs & T==`Tthree & phi2)
			 | (OP==`BCS_rel & T==`Tzero & phi1)
			 | (OP==`BCS_rel & T==`Tzero & phi2)
			 | (OP==`BCS_rel & T==`Ttwo & phi1)
			 | (OP==`BCS_rel & T==`Ttwo & phi2)
			 | (OP==`BCS_rel & T==`Tthree & phi1)
			 | (OP==`BCS_rel & T==`Tthree & phi2)
			 | (OP==`BCS_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BCS_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BCS_rel & T==`T1BranchCross & phi1)
			 | (OP==`BCS_rel & T==`T1BranchCross & phi2)
			 | (OP==`BCS_rel & T==`T1NoBranch & phi1)
			 | (OP==`BCS_rel & T==`T1NoBranch & phi2)
			 | (OP==`LDA_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDA_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`LDA_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`LDA_izy & T==`TzeroCrossPg & phi2)
			 | (OP==`LDA_izy & T==`Tone & phi1)
			 | (OP==`LDA_izy & T==`Tone & phi2)
			 | (OP==`LDA_izy & T==`Ttwo & phi1)
			 | (OP==`LDA_izy & T==`Ttwo & phi2)
			 | (OP==`LDA_izy & T==`Tthree & phi1)
			 | (OP==`LDA_izy & T==`Tthree & phi2)
			 | (OP==`LDA_izy & T==`Tfour & phi1)
			 | (OP==`LDA_izy & T==`Tfour & phi2)
			 | (OP==`LDA_izy & T==`Tfive & phi1)
			 | (OP==`LDA_izy & T==`Tfive & phi2)
			 | (OP==`LDY_zpx & T==`Tzero & phi1)
			 | (OP==`LDY_zpx & T==`Tzero & phi2)
			 | (OP==`LDY_zpx & T==`Tone & phi1)
			 | (OP==`LDY_zpx & T==`Tone & phi2)
			 | (OP==`LDY_zpx & T==`Ttwo & phi1)
			 | (OP==`LDY_zpx & T==`Ttwo & phi2)
			 | (OP==`LDY_zpx & T==`Tthree & phi1)
			 | (OP==`LDY_zpx & T==`Tthree & phi2)
			 | (OP==`LDA_zpx & T==`Tzero & phi1)
			 | (OP==`LDA_zpx & T==`Tzero & phi2)
			 | (OP==`LDA_zpx & T==`Tone & phi1)
			 | (OP==`LDA_zpx & T==`Tone & phi2)
			 | (OP==`LDA_zpx & T==`Ttwo & phi1)
			 | (OP==`LDA_zpx & T==`Ttwo & phi2)
			 | (OP==`LDA_zpx & T==`Tthree & phi1)
			 | (OP==`LDA_zpx & T==`Tthree & phi2)
			 | (OP==`LDX_zpy & T==`Tzero & phi1)
			 | (OP==`LDX_zpy & T==`Tzero & phi2)
			 | (OP==`LDX_zpy & T==`Tone & phi1)
			 | (OP==`LDX_zpy & T==`Tone & phi2)
			 | (OP==`LDX_zpy & T==`Ttwo & phi1)
			 | (OP==`LDX_zpy & T==`Ttwo & phi2)
			 | (OP==`LDX_zpy & T==`Tthree & phi1)
			 | (OP==`LDX_zpy & T==`Tthree & phi2)
			 | (OP==`CLV & T==`Tone & phi1)
			 | (OP==`CLV & T==`Tone & phi2)
			 | (OP==`CLV & T==`Ttwo & phi1)
			 | (OP==`CLV & T==`Ttwo & phi2)
			 | (OP==`LDA_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDA_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`LDA_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`LDA_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`LDA_aby & T==`Tone & phi1)
			 | (OP==`LDA_aby & T==`Tone & phi2)
			 | (OP==`LDA_aby & T==`Ttwo & phi1)
			 | (OP==`LDA_aby & T==`Ttwo & phi2)
			 | (OP==`LDA_aby & T==`Tthree & phi1)
			 | (OP==`LDA_aby & T==`Tthree & phi2)
			 | (OP==`LDA_aby & T==`Tfour & phi1)
			 | (OP==`LDA_aby & T==`Tfour & phi2)
			 | (OP==`TSX & T==`Tone & phi1)
			 | (OP==`TSX & T==`Tone & phi2)
			 | (OP==`TSX & T==`Ttwo & phi1)
			 | (OP==`TSX & T==`Ttwo & phi2)
			 | (OP==`LDY_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDY_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`LDY_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`LDY_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`LDY_abx & T==`Tone & phi1)
			 | (OP==`LDY_abx & T==`Tone & phi2)
			 | (OP==`LDY_abx & T==`Ttwo & phi1)
			 | (OP==`LDY_abx & T==`Ttwo & phi2)
			 | (OP==`LDY_abx & T==`Tthree & phi1)
			 | (OP==`LDY_abx & T==`Tthree & phi2)
			 | (OP==`LDY_abx & T==`Tfour & phi1)
			 | (OP==`LDY_abx & T==`Tfour & phi2)
			 | (OP==`LDA_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDA_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`LDA_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`LDA_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`LDA_abx & T==`Tone & phi1)
			 | (OP==`LDA_abx & T==`Tone & phi2)
			 | (OP==`LDA_abx & T==`Ttwo & phi1)
			 | (OP==`LDA_abx & T==`Ttwo & phi2)
			 | (OP==`LDA_abx & T==`Tthree & phi1)
			 | (OP==`LDA_abx & T==`Tthree & phi2)
			 | (OP==`LDA_abx & T==`Tfour & phi1)
			 | (OP==`LDA_abx & T==`Tfour & phi2)
			 | (OP==`LDX_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDX_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`LDX_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`LDX_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`LDX_aby & T==`Tone & phi1)
			 | (OP==`LDX_aby & T==`Tone & phi2)
			 | (OP==`LDX_aby & T==`Ttwo & phi1)
			 | (OP==`LDX_aby & T==`Ttwo & phi2)
			 | (OP==`LDX_aby & T==`Tthree & phi1)
			 | (OP==`LDX_aby & T==`Tthree & phi2)
			 | (OP==`LDX_aby & T==`Tfour & phi1)
			 | (OP==`LDX_aby & T==`Tfour & phi2)
			 | (OP==`CPY_imm & T==`Tone & phi1)
			 | (OP==`CPY_imm & T==`Tone & phi2)
			 | (OP==`CPY_imm & T==`Ttwo & phi1)
			 | (OP==`CPY_imm & T==`Ttwo & phi2)
			 | (OP==`CMP_izx & T==`Tzero & phi1)
			 | (OP==`CMP_izx & T==`Tzero & phi2)
			 | (OP==`CMP_izx & T==`Tone & phi1)
			 | (OP==`CMP_izx & T==`Tone & phi2)
			 | (OP==`CMP_izx & T==`Ttwo & phi1)
			 | (OP==`CMP_izx & T==`Ttwo & phi2)
			 | (OP==`CMP_izx & T==`Tthree & phi1)
			 | (OP==`CMP_izx & T==`Tthree & phi2)
			 | (OP==`CMP_izx & T==`Tfour & phi1)
			 | (OP==`CMP_izx & T==`Tfour & phi2)
			 | (OP==`CMP_izx & T==`Tfive & phi1)
			 | (OP==`CMP_izx & T==`Tfive & phi2)
			 | (OP==`CPY_zp & T==`Tzero & phi1)
			 | (OP==`CPY_zp & T==`Tzero & phi2)
			 | (OP==`CPY_zp & T==`Tone & phi1)
			 | (OP==`CPY_zp & T==`Tone & phi2)
			 | (OP==`CPY_zp & T==`Ttwo & phi1)
			 | (OP==`CPY_zp & T==`Ttwo & phi2)
			 | (OP==`CMP_zp & T==`Tzero & phi1)
			 | (OP==`CMP_zp & T==`Tzero & phi2)
			 | (OP==`CMP_zp & T==`Tone & phi1)
			 | (OP==`CMP_zp & T==`Tone & phi2)
			 | (OP==`CMP_zp & T==`Ttwo & phi1)
			 | (OP==`CMP_zp & T==`Ttwo & phi2)
			 | (OP==`DEC_zp & T==`Tzero & phi1)
			 | (OP==`DEC_zp & T==`Tzero & phi2)
			 | (OP==`DEC_zp & T==`Tone & phi1)
			 | (OP==`DEC_zp & T==`Tone & phi2)
			 | (OP==`DEC_zp & T==`Ttwo & phi1)
			 | (OP==`DEC_zp & T==`Ttwo & phi2)
			 | (OP==`DEC_zp & T==`Tthree & phi1)
			 | (OP==`DEC_zp & T==`Tthree & phi2)
			 | (OP==`DEC_zp & T==`Tfour & phi1)
			 | (OP==`DEC_zp & T==`Tfour & phi2)
			 | (OP==`INY & T==`Tone & phi1)
			 | (OP==`INY & T==`Tone & phi2)
			 | (OP==`INY & T==`Ttwo & phi1)
			 | (OP==`INY & T==`Ttwo & phi2)
			 | (OP==`CMP_imm & T==`Tone & phi1)
			 | (OP==`CMP_imm & T==`Tone & phi2)
			 | (OP==`CMP_imm & T==`Ttwo & phi1)
			 | (OP==`CMP_imm & T==`Ttwo & phi2)
			 | (OP==`DEX & T==`Tone & phi1)
			 | (OP==`DEX & T==`Tone & phi2)
			 | (OP==`DEX & T==`Ttwo & phi1)
			 | (OP==`DEX & T==`Ttwo & phi2)
			 | (OP==`CPY_abs & T==`Tzero & phi1)
			 | (OP==`CPY_abs & T==`Tzero & phi2)
			 | (OP==`CPY_abs & T==`Tone & phi1)
			 | (OP==`CPY_abs & T==`Tone & phi2)
			 | (OP==`CPY_abs & T==`Ttwo & phi1)
			 | (OP==`CPY_abs & T==`Ttwo & phi2)
			 | (OP==`CPY_abs & T==`Tthree & phi1)
			 | (OP==`CPY_abs & T==`Tthree & phi2)
			 | (OP==`CMP_abs & T==`Tzero & phi1)
			 | (OP==`CMP_abs & T==`Tzero & phi2)
			 | (OP==`CMP_abs & T==`Tone & phi1)
			 | (OP==`CMP_abs & T==`Tone & phi2)
			 | (OP==`CMP_abs & T==`Ttwo & phi1)
			 | (OP==`CMP_abs & T==`Ttwo & phi2)
			 | (OP==`CMP_abs & T==`Tthree & phi1)
			 | (OP==`CMP_abs & T==`Tthree & phi2)
			 | (OP==`DEC_abs & T==`Tzero & phi1)
			 | (OP==`DEC_abs & T==`Tzero & phi2)
			 | (OP==`DEC_abs & T==`Tone & phi1)
			 | (OP==`DEC_abs & T==`Tone & phi2)
			 | (OP==`DEC_abs & T==`Ttwo & phi1)
			 | (OP==`DEC_abs & T==`Ttwo & phi2)
			 | (OP==`DEC_abs & T==`Tthree & phi1)
			 | (OP==`DEC_abs & T==`Tthree & phi2)
			 | (OP==`DEC_abs & T==`Tfour & phi1)
			 | (OP==`DEC_abs & T==`Tfour & phi2)
			 | (OP==`DEC_abs & T==`Tfive & phi1)
			 | (OP==`DEC_abs & T==`Tfive & phi2)
			 | (OP==`BNE_rel & T==`Tzero & phi1)
			 | (OP==`BNE_rel & T==`Tzero & phi2)
			 | (OP==`BNE_rel & T==`Ttwo & phi1)
			 | (OP==`BNE_rel & T==`Ttwo & phi2)
			 | (OP==`BNE_rel & T==`Tthree & phi1)
			 | (OP==`BNE_rel & T==`Tthree & phi2)
			 | (OP==`BNE_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BNE_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BNE_rel & T==`T1BranchCross & phi1)
			 | (OP==`BNE_rel & T==`T1BranchCross & phi2)
			 | (OP==`BNE_rel & T==`T1NoBranch & phi1)
			 | (OP==`BNE_rel & T==`T1NoBranch & phi2)
			 | (OP==`CMP_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`CMP_izy & T==`TzeroCrossPg & phi2)
			 | (OP==`CMP_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`CMP_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`CMP_izy & T==`Tone & phi1)
			 | (OP==`CMP_izy & T==`Tone & phi2)
			 | (OP==`CMP_izy & T==`Ttwo & phi1)
			 | (OP==`CMP_izy & T==`Ttwo & phi2)
			 | (OP==`CMP_izy & T==`Tthree & phi1)
			 | (OP==`CMP_izy & T==`Tthree & phi2)
			 | (OP==`CMP_izy & T==`Tfour & phi1)
			 | (OP==`CMP_izy & T==`Tfour & phi2)
			 | (OP==`CMP_izy & T==`Tfive & phi1)
			 | (OP==`CMP_izy & T==`Tfive & phi2)
			 | (OP==`CMP_zpx & T==`Tzero & phi1)
			 | (OP==`CMP_zpx & T==`Tzero & phi2)
			 | (OP==`CMP_zpx & T==`Tone & phi1)
			 | (OP==`CMP_zpx & T==`Tone & phi2)
			 | (OP==`CMP_zpx & T==`Ttwo & phi1)
			 | (OP==`CMP_zpx & T==`Ttwo & phi2)
			 | (OP==`CMP_zpx & T==`Tthree & phi1)
			 | (OP==`CMP_zpx & T==`Tthree & phi2)
			 | (OP==`DEC_zpx & T==`Tzero & phi1)
			 | (OP==`DEC_zpx & T==`Tzero & phi2)
			 | (OP==`DEC_zpx & T==`Tone & phi1)
			 | (OP==`DEC_zpx & T==`Tone & phi2)
			 | (OP==`DEC_zpx & T==`Ttwo & phi1)
			 | (OP==`DEC_zpx & T==`Ttwo & phi2)
			 | (OP==`DEC_zpx & T==`Tthree & phi1)
			 | (OP==`DEC_zpx & T==`Tthree & phi2)
			 | (OP==`DEC_zpx & T==`Tfour & phi1)
			 | (OP==`DEC_zpx & T==`Tfour & phi2)
			 | (OP==`DEC_zpx & T==`Tfive & phi1)
			 | (OP==`DEC_zpx & T==`Tfive & phi2)
			 | (OP==`CLD & T==`Tone & phi1)
			 | (OP==`CLD & T==`Tone & phi2)
			 | (OP==`CLD & T==`Ttwo & phi1)
			 | (OP==`CLD & T==`Ttwo & phi2)
			 | (OP==`CMP_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`CMP_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`CMP_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`CMP_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`CMP_aby & T==`Tone & phi1)
			 | (OP==`CMP_aby & T==`Tone & phi2)
			 | (OP==`CMP_aby & T==`Ttwo & phi1)
			 | (OP==`CMP_aby & T==`Ttwo & phi2)
			 | (OP==`CMP_aby & T==`Tthree & phi1)
			 | (OP==`CMP_aby & T==`Tthree & phi2)
			 | (OP==`CMP_aby & T==`Tfour & phi1)
			 | (OP==`CMP_aby & T==`Tfour & phi2)
			 | (OP==`CMP_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`CMP_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`CMP_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`CMP_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`CMP_abx & T==`Tone & phi1)
			 | (OP==`CMP_abx & T==`Tone & phi2)
			 | (OP==`CMP_abx & T==`Ttwo & phi1)
			 | (OP==`CMP_abx & T==`Ttwo & phi2)
			 | (OP==`CMP_abx & T==`Tthree & phi1)
			 | (OP==`CMP_abx & T==`Tthree & phi2)
			 | (OP==`CMP_abx & T==`Tfour & phi1)
			 | (OP==`CMP_abx & T==`Tfour & phi2)
			 | (OP==`DEC_abx & T==`Tzero & phi1)
			 | (OP==`DEC_abx & T==`Tzero & phi2)
			 | (OP==`DEC_abx & T==`Tone & phi1)
			 | (OP==`DEC_abx & T==`Tone & phi2)
			 | (OP==`DEC_abx & T==`Ttwo & phi1)
			 | (OP==`DEC_abx & T==`Ttwo & phi2)
			 | (OP==`DEC_abx & T==`Tthree & phi1)
			 | (OP==`DEC_abx & T==`Tthree & phi2)
			 | (OP==`DEC_abx & T==`Tfour & phi1)
			 | (OP==`DEC_abx & T==`Tfour & phi2)
			 | (OP==`DEC_abx & T==`Tfive & phi1)
			 | (OP==`DEC_abx & T==`Tfive & phi2)
			 | (OP==`DEC_abx & T==`Tsix & phi1)
			 | (OP==`DEC_abx & T==`Tsix & phi2)
			 | (OP==`CPX_imm & T==`Tone & phi1)
			 | (OP==`CPX_imm & T==`Tone & phi2)
			 | (OP==`CPX_imm & T==`Ttwo & phi1)
			 | (OP==`CPX_imm & T==`Ttwo & phi2)
			 | (OP==`SBC_izx & T==`Tzero & phi1)
			 | (OP==`SBC_izx & T==`Tzero & phi2)
			 | (OP==`SBC_izx & T==`Tone & phi1)
			 | (OP==`SBC_izx & T==`Tone & phi2)
			 | (OP==`SBC_izx & T==`Ttwo & phi1)
			 | (OP==`SBC_izx & T==`Ttwo & phi2)
			 | (OP==`SBC_izx & T==`Tthree & phi1)
			 | (OP==`SBC_izx & T==`Tthree & phi2)
			 | (OP==`SBC_izx & T==`Tfour & phi1)
			 | (OP==`SBC_izx & T==`Tfour & phi2)
			 | (OP==`SBC_izx & T==`Tfive & phi1)
			 | (OP==`SBC_izx & T==`Tfive & phi2)
			 | (OP==`CPX_zp & T==`Tzero & phi1)
			 | (OP==`CPX_zp & T==`Tzero & phi2)
			 | (OP==`CPX_zp & T==`Tone & phi1)
			 | (OP==`CPX_zp & T==`Tone & phi2)
			 | (OP==`CPX_zp & T==`Ttwo & phi1)
			 | (OP==`CPX_zp & T==`Ttwo & phi2)
			 | (OP==`SBC_zp & T==`Tzero & phi1)
			 | (OP==`SBC_zp & T==`Tzero & phi2)
			 | (OP==`SBC_zp & T==`Tone & phi1)
			 | (OP==`SBC_zp & T==`Tone & phi2)
			 | (OP==`SBC_zp & T==`Ttwo & phi1)
			 | (OP==`SBC_zp & T==`Ttwo & phi2)
			 | (OP==`INC_zp & T==`Tzero & phi1)
			 | (OP==`INC_zp & T==`Tzero & phi2)
			 | (OP==`INC_zp & T==`Tone & phi1)
			 | (OP==`INC_zp & T==`Tone & phi2)
			 | (OP==`INC_zp & T==`Ttwo & phi1)
			 | (OP==`INC_zp & T==`Ttwo & phi2)
			 | (OP==`INC_zp & T==`Tthree & phi1)
			 | (OP==`INC_zp & T==`Tthree & phi2)
			 | (OP==`INC_zp & T==`Tfour & phi1)
			 | (OP==`INC_zp & T==`Tfour & phi2)
			 | (OP==`INX & T==`Tone & phi1)
			 | (OP==`INX & T==`Tone & phi2)
			 | (OP==`INX & T==`Ttwo & phi1)
			 | (OP==`INX & T==`Ttwo & phi2)
			 | (OP==`SBC_imm & T==`Tone & phi1)
			 | (OP==`SBC_imm & T==`Tone & phi2)
			 | (OP==`SBC_imm & T==`Ttwo & phi1)
			 | (OP==`SBC_imm & T==`Ttwo & phi2)
			 | (OP==`NOP & T==`Tone & phi1)
			 | (OP==`NOP & T==`Tone & phi2)
			 | (OP==`NOP & T==`Ttwo & phi1)
			 | (OP==`NOP & T==`Ttwo & phi2)
			 | (OP==`CPX_abs & T==`Tzero & phi1)
			 | (OP==`CPX_abs & T==`Tzero & phi2)
			 | (OP==`CPX_abs & T==`Tone & phi1)
			 | (OP==`CPX_abs & T==`Tone & phi2)
			 | (OP==`CPX_abs & T==`Ttwo & phi1)
			 | (OP==`CPX_abs & T==`Ttwo & phi2)
			 | (OP==`CPX_abs & T==`Tthree & phi1)
			 | (OP==`CPX_abs & T==`Tthree & phi2)
			 | (OP==`SBC_abs & T==`Tzero & phi1)
			 | (OP==`SBC_abs & T==`Tzero & phi2)
			 | (OP==`SBC_abs & T==`Tone & phi1)
			 | (OP==`SBC_abs & T==`Tone & phi2)
			 | (OP==`SBC_abs & T==`Ttwo & phi1)
			 | (OP==`SBC_abs & T==`Ttwo & phi2)
			 | (OP==`SBC_abs & T==`Tthree & phi1)
			 | (OP==`SBC_abs & T==`Tthree & phi2)
			 | (OP==`INC_abs & T==`Tzero & phi1)
			 | (OP==`INC_abs & T==`Tzero & phi2)
			 | (OP==`INC_abs & T==`Tone & phi1)
			 | (OP==`INC_abs & T==`Tone & phi2)
			 | (OP==`INC_abs & T==`Ttwo & phi1)
			 | (OP==`INC_abs & T==`Ttwo & phi2)
			 | (OP==`INC_abs & T==`Tthree & phi1)
			 | (OP==`INC_abs & T==`Tthree & phi2)
			 | (OP==`INC_abs & T==`Tfour & phi1)
			 | (OP==`INC_abs & T==`Tfour & phi2)
			 | (OP==`INC_abs & T==`Tfive & phi1)
			 | (OP==`INC_abs & T==`Tfive & phi2)
			 | (OP==`BEQ_rel & T==`Tzero & phi1)
			 | (OP==`BEQ_rel & T==`Tzero & phi2)
			 | (OP==`BEQ_rel & T==`Ttwo & phi1)
			 | (OP==`BEQ_rel & T==`Ttwo & phi2)
			 | (OP==`BEQ_rel & T==`Tthree & phi1)
			 | (OP==`BEQ_rel & T==`Tthree & phi2)
			 | (OP==`BEQ_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BEQ_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BEQ_rel & T==`T1BranchCross & phi1)
			 | (OP==`BEQ_rel & T==`T1BranchCross & phi2)
			 | (OP==`BEQ_rel & T==`T1NoBranch & phi1)
			 | (OP==`BEQ_rel & T==`T1NoBranch & phi2)
			 | (OP==`SBC_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`SBC_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`SBC_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`SBC_izy & T==`TzeroCrossPg & phi2)
			 | (OP==`SBC_izy & T==`Tone & phi1)
			 | (OP==`SBC_izy & T==`Tone & phi2)
			 | (OP==`SBC_izy & T==`Ttwo & phi1)
			 | (OP==`SBC_izy & T==`Ttwo & phi2)
			 | (OP==`SBC_izy & T==`Tthree & phi1)
			 | (OP==`SBC_izy & T==`Tthree & phi2)
			 | (OP==`SBC_izy & T==`Tfour & phi1)
			 | (OP==`SBC_izy & T==`Tfour & phi2)
			 | (OP==`SBC_izy & T==`Tfive & phi1)
			 | (OP==`SBC_izy & T==`Tfive & phi2)
			 | (OP==`SBC_zpx & T==`Tzero & phi1)
			 | (OP==`SBC_zpx & T==`Tzero & phi2)
			 | (OP==`SBC_zpx & T==`Tone & phi1)
			 | (OP==`SBC_zpx & T==`Tone & phi2)
			 | (OP==`SBC_zpx & T==`Ttwo & phi1)
			 | (OP==`SBC_zpx & T==`Ttwo & phi2)
			 | (OP==`SBC_zpx & T==`Tthree & phi1)
			 | (OP==`SBC_zpx & T==`Tthree & phi2)
			 | (OP==`INC_zpx & T==`Tzero & phi1)
			 | (OP==`INC_zpx & T==`Tzero & phi2)
			 | (OP==`INC_zpx & T==`Tone & phi1)
			 | (OP==`INC_zpx & T==`Tone & phi2)
			 | (OP==`INC_zpx & T==`Ttwo & phi1)
			 | (OP==`INC_zpx & T==`Ttwo & phi2)
			 | (OP==`INC_zpx & T==`Tthree & phi1)
			 | (OP==`INC_zpx & T==`Tthree & phi2)
			 | (OP==`INC_zpx & T==`Tfour & phi1)
			 | (OP==`INC_zpx & T==`Tfour & phi2)
			 | (OP==`INC_zpx & T==`Tfive & phi1)
			 | (OP==`INC_zpx & T==`Tfive & phi2)
			 | (OP==`SED & T==`Tone & phi1)
			 | (OP==`SED & T==`Tone & phi2)
			 | (OP==`SED & T==`Ttwo & phi1)
			 | (OP==`SED & T==`Ttwo & phi2)
			 | (OP==`SBC_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`SBC_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`SBC_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`SBC_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`SBC_aby & T==`Tone & phi1)
			 | (OP==`SBC_aby & T==`Tone & phi2)
			 | (OP==`SBC_aby & T==`Ttwo & phi1)
			 | (OP==`SBC_aby & T==`Ttwo & phi2)
			 | (OP==`SBC_aby & T==`Tthree & phi1)
			 | (OP==`SBC_aby & T==`Tthree & phi2)
			 | (OP==`SBC_aby & T==`Tfour & phi1)
			 | (OP==`SBC_aby & T==`Tfour & phi2)
			 | (OP==`SBC_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`SBC_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`SBC_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`SBC_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`SBC_abx & T==`Tone & phi1)
			 | (OP==`SBC_abx & T==`Tone & phi2)
			 | (OP==`SBC_abx & T==`Ttwo & phi1)
			 | (OP==`SBC_abx & T==`Ttwo & phi2)
			 | (OP==`SBC_abx & T==`Tthree & phi1)
			 | (OP==`SBC_abx & T==`Tthree & phi2)
			 | (OP==`SBC_abx & T==`Tfour & phi1)
			 | (OP==`SBC_abx & T==`Tfour & phi2)
			 | (OP==`INC_abx & T==`Tzero & phi1)
			 | (OP==`INC_abx & T==`Tzero & phi2)
			 | (OP==`INC_abx & T==`Tone & phi1)
			 | (OP==`INC_abx & T==`Tone & phi2)
			 | (OP==`INC_abx & T==`Ttwo & phi1)
			 | (OP==`INC_abx & T==`Ttwo & phi2)
			 | (OP==`INC_abx & T==`Tthree & phi1)
			 | (OP==`INC_abx & T==`Tthree & phi2)
			 | (OP==`INC_abx & T==`Tfour & phi1)
			 | (OP==`INC_abx & T==`Tfour & phi2)
			 | (OP==`INC_abx & T==`Tfive & phi1)
			 | (OP==`INC_abx & T==`Tfive & phi2)
			 | (OP==`INC_abx & T==`Tsix & phi1)
			 | (OP==`INC_abx & T==`Tsix & phi2)
			;

assign control[`nDSA] = (OP==`BRK & T==`Tzero & phi1)
			 | (OP==`BRK & T==`Tzero & phi2)
			 | (OP==`BRK & T==`Tone & phi1)
			 | (OP==`BRK & T==`Tone & phi2)
			 | (OP==`BRK & T==`Ttwo & phi1)
			 | (OP==`BRK & T==`Ttwo & phi2)
			 | (OP==`BRK & T==`Tthree & phi1)
			 | (OP==`BRK & T==`Tthree & phi2)
			 | (OP==`BRK & T==`Tfour & phi1)
			 | (OP==`BRK & T==`Tfour & phi2)
			 | (OP==`BRK & T==`Tfive & phi1)
			 | (OP==`BRK & T==`Tfive & phi2)
			 | (OP==`BRK & T==`Tsix & phi1)
			 | (OP==`BRK & T==`Tsix & phi2)
			 | (OP==`ORA_izx & T==`Tzero & phi1)
			 | (OP==`ORA_izx & T==`Tzero & phi2)
			 | (OP==`ORA_izx & T==`Tone & phi1)
			 | (OP==`ORA_izx & T==`Tone & phi2)
			 | (OP==`ORA_izx & T==`Ttwo & phi1)
			 | (OP==`ORA_izx & T==`Ttwo & phi2)
			 | (OP==`ORA_izx & T==`Tthree & phi1)
			 | (OP==`ORA_izx & T==`Tthree & phi2)
			 | (OP==`ORA_izx & T==`Tfour & phi1)
			 | (OP==`ORA_izx & T==`Tfour & phi2)
			 | (OP==`ORA_izx & T==`Tfive & phi1)
			 | (OP==`ORA_izx & T==`Tfive & phi2)
			 | (OP==`ORA_zp & T==`Tzero & phi1)
			 | (OP==`ORA_zp & T==`Tzero & phi2)
			 | (OP==`ORA_zp & T==`Tone & phi1)
			 | (OP==`ORA_zp & T==`Tone & phi2)
			 | (OP==`ORA_zp & T==`Ttwo & phi1)
			 | (OP==`ORA_zp & T==`Ttwo & phi2)
			 | (OP==`ASL_zp & T==`Tzero & phi1)
			 | (OP==`ASL_zp & T==`Tzero & phi2)
			 | (OP==`ASL_zp & T==`Tone & phi1)
			 | (OP==`ASL_zp & T==`Tone & phi2)
			 | (OP==`ASL_zp & T==`Ttwo & phi1)
			 | (OP==`ASL_zp & T==`Ttwo & phi2)
			 | (OP==`ASL_zp & T==`Tthree & phi1)
			 | (OP==`ASL_zp & T==`Tthree & phi2)
			 | (OP==`ASL_zp & T==`Tfour & phi1)
			 | (OP==`ASL_zp & T==`Tfour & phi2)
			 | (OP==`PHP & T==`Tzero & phi1)
			 | (OP==`PHP & T==`Tzero & phi2)
			 | (OP==`PHP & T==`Tone & phi1)
			 | (OP==`PHP & T==`Tone & phi2)
			 | (OP==`PHP & T==`Ttwo & phi1)
			 | (OP==`PHP & T==`Ttwo & phi2)
			 | (OP==`ORA_imm & T==`Tone & phi1)
			 | (OP==`ORA_imm & T==`Tone & phi2)
			 | (OP==`ORA_imm & T==`Ttwo & phi1)
			 | (OP==`ORA_imm & T==`Ttwo & phi2)
			 | (OP==`ASL & T==`Tone & phi1)
			 | (OP==`ASL & T==`Tone & phi2)
			 | (OP==`ASL & T==`Ttwo & phi1)
			 | (OP==`ASL & T==`Ttwo & phi2)
			 | (OP==`ORA_abs & T==`Tzero & phi1)
			 | (OP==`ORA_abs & T==`Tzero & phi2)
			 | (OP==`ORA_abs & T==`Tone & phi1)
			 | (OP==`ORA_abs & T==`Tone & phi2)
			 | (OP==`ORA_abs & T==`Ttwo & phi1)
			 | (OP==`ORA_abs & T==`Ttwo & phi2)
			 | (OP==`ORA_abs & T==`Tthree & phi1)
			 | (OP==`ORA_abs & T==`Tthree & phi2)
			 | (OP==`ASL_abs & T==`Tzero & phi1)
			 | (OP==`ASL_abs & T==`Tzero & phi2)
			 | (OP==`ASL_abs & T==`Tone & phi1)
			 | (OP==`ASL_abs & T==`Tone & phi2)
			 | (OP==`ASL_abs & T==`Ttwo & phi1)
			 | (OP==`ASL_abs & T==`Ttwo & phi2)
			 | (OP==`ASL_abs & T==`Tthree & phi1)
			 | (OP==`ASL_abs & T==`Tthree & phi2)
			 | (OP==`ASL_abs & T==`Tfour & phi1)
			 | (OP==`ASL_abs & T==`Tfour & phi2)
			 | (OP==`ASL_abs & T==`Tfive & phi1)
			 | (OP==`ASL_abs & T==`Tfive & phi2)
			 | (OP==`BPL_rel & T==`Tzero & phi1)
			 | (OP==`BPL_rel & T==`Tzero & phi2)
			 | (OP==`BPL_rel & T==`Ttwo & phi1)
			 | (OP==`BPL_rel & T==`Ttwo & phi2)
			 | (OP==`BPL_rel & T==`Tthree & phi1)
			 | (OP==`BPL_rel & T==`Tthree & phi2)
			 | (OP==`BPL_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BPL_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BPL_rel & T==`T1BranchCross & phi1)
			 | (OP==`BPL_rel & T==`T1BranchCross & phi2)
			 | (OP==`BPL_rel & T==`T1NoBranch & phi1)
			 | (OP==`BPL_rel & T==`T1NoBranch & phi2)
			 | (OP==`ORA_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`ORA_izy & T==`TzeroCrossPg & phi2)
			 | (OP==`ORA_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ORA_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`ORA_izy & T==`Tone & phi1)
			 | (OP==`ORA_izy & T==`Tone & phi2)
			 | (OP==`ORA_izy & T==`Ttwo & phi1)
			 | (OP==`ORA_izy & T==`Ttwo & phi2)
			 | (OP==`ORA_izy & T==`Tthree & phi1)
			 | (OP==`ORA_izy & T==`Tthree & phi2)
			 | (OP==`ORA_izy & T==`Tfour & phi1)
			 | (OP==`ORA_izy & T==`Tfour & phi2)
			 | (OP==`ORA_izy & T==`Tfive & phi1)
			 | (OP==`ORA_izy & T==`Tfive & phi2)
			 | (OP==`ORA_zpx & T==`Tzero & phi1)
			 | (OP==`ORA_zpx & T==`Tzero & phi2)
			 | (OP==`ORA_zpx & T==`Tone & phi1)
			 | (OP==`ORA_zpx & T==`Tone & phi2)
			 | (OP==`ORA_zpx & T==`Ttwo & phi1)
			 | (OP==`ORA_zpx & T==`Ttwo & phi2)
			 | (OP==`ORA_zpx & T==`Tthree & phi1)
			 | (OP==`ORA_zpx & T==`Tthree & phi2)
			 | (OP==`ASL_zpx & T==`Tzero & phi1)
			 | (OP==`ASL_zpx & T==`Tzero & phi2)
			 | (OP==`ASL_zpx & T==`Tone & phi1)
			 | (OP==`ASL_zpx & T==`Tone & phi2)
			 | (OP==`ASL_zpx & T==`Ttwo & phi1)
			 | (OP==`ASL_zpx & T==`Ttwo & phi2)
			 | (OP==`ASL_zpx & T==`Tthree & phi1)
			 | (OP==`ASL_zpx & T==`Tthree & phi2)
			 | (OP==`ASL_zpx & T==`Tfour & phi1)
			 | (OP==`ASL_zpx & T==`Tfour & phi2)
			 | (OP==`ASL_zpx & T==`Tfive & phi1)
			 | (OP==`ASL_zpx & T==`Tfive & phi2)
			 | (OP==`CLC & T==`Tone & phi1)
			 | (OP==`CLC & T==`Tone & phi2)
			 | (OP==`CLC & T==`Ttwo & phi1)
			 | (OP==`CLC & T==`Ttwo & phi2)
			 | (OP==`ORA_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ORA_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`ORA_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`ORA_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`ORA_aby & T==`Tone & phi1)
			 | (OP==`ORA_aby & T==`Tone & phi2)
			 | (OP==`ORA_aby & T==`Ttwo & phi1)
			 | (OP==`ORA_aby & T==`Ttwo & phi2)
			 | (OP==`ORA_aby & T==`Tthree & phi1)
			 | (OP==`ORA_aby & T==`Tthree & phi2)
			 | (OP==`ORA_aby & T==`Tfour & phi1)
			 | (OP==`ORA_aby & T==`Tfour & phi2)
			 | (OP==`ORA_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ORA_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`ORA_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`ORA_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`ORA_abx & T==`Tone & phi1)
			 | (OP==`ORA_abx & T==`Tone & phi2)
			 | (OP==`ORA_abx & T==`Ttwo & phi1)
			 | (OP==`ORA_abx & T==`Ttwo & phi2)
			 | (OP==`ORA_abx & T==`Tthree & phi1)
			 | (OP==`ORA_abx & T==`Tthree & phi2)
			 | (OP==`ORA_abx & T==`Tfour & phi1)
			 | (OP==`ORA_abx & T==`Tfour & phi2)
			 | (OP==`ASL_abx & T==`Tzero & phi1)
			 | (OP==`ASL_abx & T==`Tzero & phi2)
			 | (OP==`ASL_abx & T==`Tone & phi1)
			 | (OP==`ASL_abx & T==`Tone & phi2)
			 | (OP==`ASL_abx & T==`Ttwo & phi1)
			 | (OP==`ASL_abx & T==`Ttwo & phi2)
			 | (OP==`ASL_abx & T==`Tthree & phi1)
			 | (OP==`ASL_abx & T==`Tthree & phi2)
			 | (OP==`ASL_abx & T==`Tfour & phi1)
			 | (OP==`ASL_abx & T==`Tfour & phi2)
			 | (OP==`ASL_abx & T==`Tfive & phi1)
			 | (OP==`ASL_abx & T==`Tfive & phi2)
			 | (OP==`ASL_abx & T==`Tsix & phi1)
			 | (OP==`ASL_abx & T==`Tsix & phi2)
			 | (OP==`JSR_abs & T==`Tzero & phi1)
			 | (OP==`JSR_abs & T==`Tzero & phi2)
			 | (OP==`JSR_abs & T==`Tone & phi1)
			 | (OP==`JSR_abs & T==`Tone & phi2)
			 | (OP==`JSR_abs & T==`Ttwo & phi1)
			 | (OP==`JSR_abs & T==`Ttwo & phi2)
			 | (OP==`JSR_abs & T==`Tthree & phi1)
			 | (OP==`JSR_abs & T==`Tthree & phi2)
			 | (OP==`JSR_abs & T==`Tfour & phi1)
			 | (OP==`JSR_abs & T==`Tfour & phi2)
			 | (OP==`JSR_abs & T==`Tfive & phi1)
			 | (OP==`JSR_abs & T==`Tfive & phi2)
			 | (OP==`AND_izx & T==`Tzero & phi1)
			 | (OP==`AND_izx & T==`Tzero & phi2)
			 | (OP==`AND_izx & T==`Tone & phi1)
			 | (OP==`AND_izx & T==`Tone & phi2)
			 | (OP==`AND_izx & T==`Ttwo & phi1)
			 | (OP==`AND_izx & T==`Ttwo & phi2)
			 | (OP==`AND_izx & T==`Tthree & phi1)
			 | (OP==`AND_izx & T==`Tthree & phi2)
			 | (OP==`AND_izx & T==`Tfour & phi1)
			 | (OP==`AND_izx & T==`Tfour & phi2)
			 | (OP==`AND_izx & T==`Tfive & phi1)
			 | (OP==`AND_izx & T==`Tfive & phi2)
			 | (OP==`BIT_zp & T==`Tzero & phi1)
			 | (OP==`BIT_zp & T==`Tzero & phi2)
			 | (OP==`BIT_zp & T==`Tone & phi1)
			 | (OP==`BIT_zp & T==`Tone & phi2)
			 | (OP==`BIT_zp & T==`Ttwo & phi1)
			 | (OP==`BIT_zp & T==`Ttwo & phi2)
			 | (OP==`AND_zp & T==`Tzero & phi1)
			 | (OP==`AND_zp & T==`Tzero & phi2)
			 | (OP==`AND_zp & T==`Tone & phi1)
			 | (OP==`AND_zp & T==`Tone & phi2)
			 | (OP==`AND_zp & T==`Ttwo & phi1)
			 | (OP==`AND_zp & T==`Ttwo & phi2)
			 | (OP==`ROL_zp & T==`Tzero & phi1)
			 | (OP==`ROL_zp & T==`Tzero & phi2)
			 | (OP==`ROL_zp & T==`Tone & phi1)
			 | (OP==`ROL_zp & T==`Tone & phi2)
			 | (OP==`ROL_zp & T==`Ttwo & phi1)
			 | (OP==`ROL_zp & T==`Ttwo & phi2)
			 | (OP==`ROL_zp & T==`Tthree & phi1)
			 | (OP==`ROL_zp & T==`Tthree & phi2)
			 | (OP==`ROL_zp & T==`Tfour & phi1)
			 | (OP==`ROL_zp & T==`Tfour & phi2)
			 | (OP==`PLP & T==`Tzero & phi1)
			 | (OP==`PLP & T==`Tzero & phi2)
			 | (OP==`PLP & T==`Tone & phi1)
			 | (OP==`PLP & T==`Tone & phi2)
			 | (OP==`PLP & T==`Ttwo & phi1)
			 | (OP==`PLP & T==`Ttwo & phi2)
			 | (OP==`PLP & T==`Tthree & phi1)
			 | (OP==`PLP & T==`Tthree & phi2)
			 | (OP==`AND_imm & T==`Tone & phi1)
			 | (OP==`AND_imm & T==`Tone & phi2)
			 | (OP==`AND_imm & T==`Ttwo & phi1)
			 | (OP==`AND_imm & T==`Ttwo & phi2)
			 | (OP==`ROL & T==`Tone & phi1)
			 | (OP==`ROL & T==`Tone & phi2)
			 | (OP==`ROL & T==`Ttwo & phi1)
			 | (OP==`ROL & T==`Ttwo & phi2)
			 | (OP==`BIT_abs & T==`Tzero & phi1)
			 | (OP==`BIT_abs & T==`Tzero & phi2)
			 | (OP==`BIT_abs & T==`Tone & phi1)
			 | (OP==`BIT_abs & T==`Tone & phi2)
			 | (OP==`BIT_abs & T==`Ttwo & phi1)
			 | (OP==`BIT_abs & T==`Ttwo & phi2)
			 | (OP==`BIT_abs & T==`Tthree & phi1)
			 | (OP==`BIT_abs & T==`Tthree & phi2)
			 | (OP==`AND_abs & T==`Tzero & phi1)
			 | (OP==`AND_abs & T==`Tzero & phi2)
			 | (OP==`AND_abs & T==`Tone & phi1)
			 | (OP==`AND_abs & T==`Tone & phi2)
			 | (OP==`AND_abs & T==`Ttwo & phi1)
			 | (OP==`AND_abs & T==`Ttwo & phi2)
			 | (OP==`AND_abs & T==`Tthree & phi1)
			 | (OP==`AND_abs & T==`Tthree & phi2)
			 | (OP==`ROL_abs & T==`Tzero & phi1)
			 | (OP==`ROL_abs & T==`Tzero & phi2)
			 | (OP==`ROL_abs & T==`Tone & phi1)
			 | (OP==`ROL_abs & T==`Tone & phi2)
			 | (OP==`ROL_abs & T==`Ttwo & phi1)
			 | (OP==`ROL_abs & T==`Ttwo & phi2)
			 | (OP==`ROL_abs & T==`Tthree & phi1)
			 | (OP==`ROL_abs & T==`Tthree & phi2)
			 | (OP==`ROL_abs & T==`Tfour & phi1)
			 | (OP==`ROL_abs & T==`Tfour & phi2)
			 | (OP==`ROL_abs & T==`Tfive & phi1)
			 | (OP==`ROL_abs & T==`Tfive & phi2)
			 | (OP==`BMI_rel & T==`Tzero & phi1)
			 | (OP==`BMI_rel & T==`Tzero & phi2)
			 | (OP==`BMI_rel & T==`Ttwo & phi1)
			 | (OP==`BMI_rel & T==`Ttwo & phi2)
			 | (OP==`BMI_rel & T==`Tthree & phi1)
			 | (OP==`BMI_rel & T==`Tthree & phi2)
			 | (OP==`BMI_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BMI_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BMI_rel & T==`T1BranchCross & phi1)
			 | (OP==`BMI_rel & T==`T1BranchCross & phi2)
			 | (OP==`BMI_rel & T==`T1NoBranch & phi1)
			 | (OP==`BMI_rel & T==`T1NoBranch & phi2)
			 | (OP==`AND_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`AND_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`AND_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`AND_izy & T==`TzeroCrossPg & phi2)
			 | (OP==`AND_izy & T==`Tone & phi1)
			 | (OP==`AND_izy & T==`Tone & phi2)
			 | (OP==`AND_izy & T==`Ttwo & phi1)
			 | (OP==`AND_izy & T==`Ttwo & phi2)
			 | (OP==`AND_izy & T==`Tthree & phi1)
			 | (OP==`AND_izy & T==`Tthree & phi2)
			 | (OP==`AND_izy & T==`Tfour & phi1)
			 | (OP==`AND_izy & T==`Tfour & phi2)
			 | (OP==`AND_izy & T==`Tfive & phi1)
			 | (OP==`AND_izy & T==`Tfive & phi2)
			 | (OP==`AND_zpx & T==`Tzero & phi1)
			 | (OP==`AND_zpx & T==`Tzero & phi2)
			 | (OP==`AND_zpx & T==`Tone & phi1)
			 | (OP==`AND_zpx & T==`Tone & phi2)
			 | (OP==`AND_zpx & T==`Ttwo & phi1)
			 | (OP==`AND_zpx & T==`Ttwo & phi2)
			 | (OP==`AND_zpx & T==`Tthree & phi1)
			 | (OP==`AND_zpx & T==`Tthree & phi2)
			 | (OP==`ROL_zpx & T==`Tzero & phi1)
			 | (OP==`ROL_zpx & T==`Tzero & phi2)
			 | (OP==`ROL_zpx & T==`Tone & phi1)
			 | (OP==`ROL_zpx & T==`Tone & phi2)
			 | (OP==`ROL_zpx & T==`Ttwo & phi1)
			 | (OP==`ROL_zpx & T==`Ttwo & phi2)
			 | (OP==`ROL_zpx & T==`Tthree & phi1)
			 | (OP==`ROL_zpx & T==`Tthree & phi2)
			 | (OP==`ROL_zpx & T==`Tfour & phi1)
			 | (OP==`ROL_zpx & T==`Tfour & phi2)
			 | (OP==`ROL_zpx & T==`Tfive & phi1)
			 | (OP==`ROL_zpx & T==`Tfive & phi2)
			 | (OP==`SEC & T==`Tone & phi1)
			 | (OP==`SEC & T==`Tone & phi2)
			 | (OP==`SEC & T==`Ttwo & phi1)
			 | (OP==`SEC & T==`Ttwo & phi2)
			 | (OP==`AND_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`AND_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`AND_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`AND_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`AND_aby & T==`Tone & phi1)
			 | (OP==`AND_aby & T==`Tone & phi2)
			 | (OP==`AND_aby & T==`Ttwo & phi1)
			 | (OP==`AND_aby & T==`Ttwo & phi2)
			 | (OP==`AND_aby & T==`Tthree & phi1)
			 | (OP==`AND_aby & T==`Tthree & phi2)
			 | (OP==`AND_aby & T==`Tfour & phi1)
			 | (OP==`AND_aby & T==`Tfour & phi2)
			 | (OP==`AND_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`AND_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`AND_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`AND_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`AND_abx & T==`Tone & phi1)
			 | (OP==`AND_abx & T==`Tone & phi2)
			 | (OP==`AND_abx & T==`Ttwo & phi1)
			 | (OP==`AND_abx & T==`Ttwo & phi2)
			 | (OP==`AND_abx & T==`Tthree & phi1)
			 | (OP==`AND_abx & T==`Tthree & phi2)
			 | (OP==`AND_abx & T==`Tfour & phi1)
			 | (OP==`AND_abx & T==`Tfour & phi2)
			 | (OP==`ROL_abx & T==`Tzero & phi1)
			 | (OP==`ROL_abx & T==`Tzero & phi2)
			 | (OP==`ROL_abx & T==`Tone & phi1)
			 | (OP==`ROL_abx & T==`Tone & phi2)
			 | (OP==`ROL_abx & T==`Ttwo & phi1)
			 | (OP==`ROL_abx & T==`Ttwo & phi2)
			 | (OP==`ROL_abx & T==`Tthree & phi1)
			 | (OP==`ROL_abx & T==`Tthree & phi2)
			 | (OP==`ROL_abx & T==`Tfour & phi1)
			 | (OP==`ROL_abx & T==`Tfour & phi2)
			 | (OP==`ROL_abx & T==`Tfive & phi1)
			 | (OP==`ROL_abx & T==`Tfive & phi2)
			 | (OP==`ROL_abx & T==`Tsix & phi1)
			 | (OP==`ROL_abx & T==`Tsix & phi2)
			 | (OP==`RTI & T==`Tzero & phi1)
			 | (OP==`RTI & T==`Tzero & phi2)
			 | (OP==`RTI & T==`Tone & phi1)
			 | (OP==`RTI & T==`Tone & phi2)
			 | (OP==`RTI & T==`Ttwo & phi1)
			 | (OP==`RTI & T==`Ttwo & phi2)
			 | (OP==`RTI & T==`Tthree & phi1)
			 | (OP==`RTI & T==`Tthree & phi2)
			 | (OP==`RTI & T==`Tfour & phi1)
			 | (OP==`RTI & T==`Tfour & phi2)
			 | (OP==`RTI & T==`Tfive & phi1)
			 | (OP==`RTI & T==`Tfive & phi2)
			 | (OP==`EOR_izx & T==`Tzero & phi1)
			 | (OP==`EOR_izx & T==`Tzero & phi2)
			 | (OP==`EOR_izx & T==`Tone & phi1)
			 | (OP==`EOR_izx & T==`Tone & phi2)
			 | (OP==`EOR_izx & T==`Ttwo & phi1)
			 | (OP==`EOR_izx & T==`Ttwo & phi2)
			 | (OP==`EOR_izx & T==`Tthree & phi1)
			 | (OP==`EOR_izx & T==`Tthree & phi2)
			 | (OP==`EOR_izx & T==`Tfour & phi1)
			 | (OP==`EOR_izx & T==`Tfour & phi2)
			 | (OP==`EOR_izx & T==`Tfive & phi1)
			 | (OP==`EOR_izx & T==`Tfive & phi2)
			 | (OP==`EOR_zp & T==`Tzero & phi1)
			 | (OP==`EOR_zp & T==`Tzero & phi2)
			 | (OP==`EOR_zp & T==`Tone & phi1)
			 | (OP==`EOR_zp & T==`Tone & phi2)
			 | (OP==`EOR_zp & T==`Ttwo & phi1)
			 | (OP==`EOR_zp & T==`Ttwo & phi2)
			 | (OP==`LSR_zp & T==`Tzero & phi1)
			 | (OP==`LSR_zp & T==`Tzero & phi2)
			 | (OP==`LSR_zp & T==`Tone & phi1)
			 | (OP==`LSR_zp & T==`Tone & phi2)
			 | (OP==`LSR_zp & T==`Ttwo & phi1)
			 | (OP==`LSR_zp & T==`Ttwo & phi2)
			 | (OP==`LSR_zp & T==`Tthree & phi1)
			 | (OP==`LSR_zp & T==`Tthree & phi2)
			 | (OP==`LSR_zp & T==`Tfour & phi1)
			 | (OP==`LSR_zp & T==`Tfour & phi2)
			 | (OP==`PHA & T==`Tzero & phi1)
			 | (OP==`PHA & T==`Tzero & phi2)
			 | (OP==`PHA & T==`Tone & phi1)
			 | (OP==`PHA & T==`Tone & phi2)
			 | (OP==`PHA & T==`Ttwo & phi1)
			 | (OP==`PHA & T==`Ttwo & phi2)
			 | (OP==`EOR_imm & T==`Tone & phi1)
			 | (OP==`EOR_imm & T==`Tone & phi2)
			 | (OP==`EOR_imm & T==`Ttwo & phi1)
			 | (OP==`EOR_imm & T==`Ttwo & phi2)
			 | (OP==`LSR & T==`Tone & phi1)
			 | (OP==`LSR & T==`Tone & phi2)
			 | (OP==`LSR & T==`Ttwo & phi1)
			 | (OP==`LSR & T==`Ttwo & phi2)
			 | (OP==`JMP_abs & T==`Tzero & phi1)
			 | (OP==`JMP_abs & T==`Tzero & phi2)
			 | (OP==`JMP_abs & T==`Tone & phi1)
			 | (OP==`JMP_abs & T==`Tone & phi2)
			 | (OP==`JMP_abs & T==`Ttwo & phi1)
			 | (OP==`JMP_abs & T==`Ttwo & phi2)
			 | (OP==`EOR_abs & T==`Tzero & phi1)
			 | (OP==`EOR_abs & T==`Tzero & phi2)
			 | (OP==`EOR_abs & T==`Tone & phi1)
			 | (OP==`EOR_abs & T==`Tone & phi2)
			 | (OP==`EOR_abs & T==`Ttwo & phi1)
			 | (OP==`EOR_abs & T==`Ttwo & phi2)
			 | (OP==`EOR_abs & T==`Tthree & phi1)
			 | (OP==`EOR_abs & T==`Tthree & phi2)
			 | (OP==`LSR_abs & T==`Tzero & phi1)
			 | (OP==`LSR_abs & T==`Tzero & phi2)
			 | (OP==`LSR_abs & T==`Tone & phi1)
			 | (OP==`LSR_abs & T==`Tone & phi2)
			 | (OP==`LSR_abs & T==`Ttwo & phi1)
			 | (OP==`LSR_abs & T==`Ttwo & phi2)
			 | (OP==`LSR_abs & T==`Tthree & phi1)
			 | (OP==`LSR_abs & T==`Tthree & phi2)
			 | (OP==`LSR_abs & T==`Tfour & phi1)
			 | (OP==`LSR_abs & T==`Tfour & phi2)
			 | (OP==`LSR_abs & T==`Tfive & phi1)
			 | (OP==`LSR_abs & T==`Tfive & phi2)
			 | (OP==`BVC_rel & T==`Tzero & phi1)
			 | (OP==`BVC_rel & T==`Tzero & phi2)
			 | (OP==`BVC_rel & T==`Ttwo & phi1)
			 | (OP==`BVC_rel & T==`Ttwo & phi2)
			 | (OP==`BVC_rel & T==`Tthree & phi1)
			 | (OP==`BVC_rel & T==`Tthree & phi2)
			 | (OP==`BVC_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BVC_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BVC_rel & T==`T1BranchCross & phi1)
			 | (OP==`BVC_rel & T==`T1BranchCross & phi2)
			 | (OP==`BVC_rel & T==`T1NoBranch & phi1)
			 | (OP==`BVC_rel & T==`T1NoBranch & phi2)
			 | (OP==`EOR_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`EOR_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`EOR_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`EOR_izy & T==`TzeroCrossPg & phi2)
			 | (OP==`EOR_izy & T==`Tone & phi1)
			 | (OP==`EOR_izy & T==`Tone & phi2)
			 | (OP==`EOR_izy & T==`Ttwo & phi1)
			 | (OP==`EOR_izy & T==`Ttwo & phi2)
			 | (OP==`EOR_izy & T==`Tthree & phi1)
			 | (OP==`EOR_izy & T==`Tthree & phi2)
			 | (OP==`EOR_izy & T==`Tfour & phi1)
			 | (OP==`EOR_izy & T==`Tfour & phi2)
			 | (OP==`EOR_izy & T==`Tfive & phi1)
			 | (OP==`EOR_izy & T==`Tfive & phi2)
			 | (OP==`EOR_zpx & T==`Tzero & phi1)
			 | (OP==`EOR_zpx & T==`Tzero & phi2)
			 | (OP==`EOR_zpx & T==`Tone & phi1)
			 | (OP==`EOR_zpx & T==`Tone & phi2)
			 | (OP==`EOR_zpx & T==`Ttwo & phi1)
			 | (OP==`EOR_zpx & T==`Ttwo & phi2)
			 | (OP==`EOR_zpx & T==`Tthree & phi1)
			 | (OP==`EOR_zpx & T==`Tthree & phi2)
			 | (OP==`LSR_zpx & T==`Tzero & phi1)
			 | (OP==`LSR_zpx & T==`Tzero & phi2)
			 | (OP==`LSR_zpx & T==`Tone & phi1)
			 | (OP==`LSR_zpx & T==`Tone & phi2)
			 | (OP==`LSR_zpx & T==`Ttwo & phi1)
			 | (OP==`LSR_zpx & T==`Ttwo & phi2)
			 | (OP==`LSR_zpx & T==`Tthree & phi1)
			 | (OP==`LSR_zpx & T==`Tthree & phi2)
			 | (OP==`LSR_zpx & T==`Tfour & phi1)
			 | (OP==`LSR_zpx & T==`Tfour & phi2)
			 | (OP==`LSR_zpx & T==`Tfive & phi1)
			 | (OP==`LSR_zpx & T==`Tfive & phi2)
			 | (OP==`CLI & T==`Tone & phi1)
			 | (OP==`CLI & T==`Tone & phi2)
			 | (OP==`CLI & T==`Ttwo & phi1)
			 | (OP==`CLI & T==`Ttwo & phi2)
			 | (OP==`EOR_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`EOR_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`EOR_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`EOR_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`EOR_aby & T==`Tone & phi1)
			 | (OP==`EOR_aby & T==`Tone & phi2)
			 | (OP==`EOR_aby & T==`Ttwo & phi1)
			 | (OP==`EOR_aby & T==`Ttwo & phi2)
			 | (OP==`EOR_aby & T==`Tthree & phi1)
			 | (OP==`EOR_aby & T==`Tthree & phi2)
			 | (OP==`EOR_aby & T==`Tfour & phi1)
			 | (OP==`EOR_aby & T==`Tfour & phi2)
			 | (OP==`EOR_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`EOR_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`EOR_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`EOR_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`EOR_abx & T==`Tone & phi1)
			 | (OP==`EOR_abx & T==`Tone & phi2)
			 | (OP==`EOR_abx & T==`Ttwo & phi1)
			 | (OP==`EOR_abx & T==`Ttwo & phi2)
			 | (OP==`EOR_abx & T==`Tthree & phi1)
			 | (OP==`EOR_abx & T==`Tthree & phi2)
			 | (OP==`EOR_abx & T==`Tfour & phi1)
			 | (OP==`EOR_abx & T==`Tfour & phi2)
			 | (OP==`LSR_abx & T==`Tzero & phi1)
			 | (OP==`LSR_abx & T==`Tzero & phi2)
			 | (OP==`LSR_abx & T==`Tone & phi1)
			 | (OP==`LSR_abx & T==`Tone & phi2)
			 | (OP==`LSR_abx & T==`Ttwo & phi1)
			 | (OP==`LSR_abx & T==`Ttwo & phi2)
			 | (OP==`LSR_abx & T==`Tthree & phi1)
			 | (OP==`LSR_abx & T==`Tthree & phi2)
			 | (OP==`LSR_abx & T==`Tfour & phi1)
			 | (OP==`LSR_abx & T==`Tfour & phi2)
			 | (OP==`LSR_abx & T==`Tfive & phi1)
			 | (OP==`LSR_abx & T==`Tfive & phi2)
			 | (OP==`LSR_abx & T==`Tsix & phi1)
			 | (OP==`LSR_abx & T==`Tsix & phi2)
			 | (OP==`RTS & T==`Tzero & phi1)
			 | (OP==`RTS & T==`Tzero & phi2)
			 | (OP==`RTS & T==`Tone & phi1)
			 | (OP==`RTS & T==`Tone & phi2)
			 | (OP==`RTS & T==`Ttwo & phi1)
			 | (OP==`RTS & T==`Ttwo & phi2)
			 | (OP==`RTS & T==`Tthree & phi1)
			 | (OP==`RTS & T==`Tthree & phi2)
			 | (OP==`RTS & T==`Tfour & phi1)
			 | (OP==`RTS & T==`Tfour & phi2)
			 | (OP==`RTS & T==`Tfive & phi1)
			 | (OP==`RTS & T==`Tfive & phi2)
			 | (OP==`ADC_izx & T==`Tzero & phi1)
			 | (OP==`ADC_izx & T==`Tzero & phi2)
			 | (OP==`ADC_izx & T==`Tone & phi1)
			 | (OP==`ADC_izx & T==`Tone & phi2)
			 | (OP==`ADC_izx & T==`Ttwo & phi1)
			 | (OP==`ADC_izx & T==`Ttwo & phi2)
			 | (OP==`ADC_izx & T==`Tthree & phi1)
			 | (OP==`ADC_izx & T==`Tthree & phi2)
			 | (OP==`ADC_izx & T==`Tfour & phi1)
			 | (OP==`ADC_izx & T==`Tfour & phi2)
			 | (OP==`ADC_izx & T==`Tfive & phi1)
			 | (OP==`ADC_izx & T==`Tfive & phi2)
			 | (OP==`ADC_zp & T==`Tzero & phi1)
			 | (OP==`ADC_zp & T==`Tzero & phi2)
			 | (OP==`ADC_zp & T==`Tone & phi1)
			 | (OP==`ADC_zp & T==`Tone & phi2)
			 | (OP==`ADC_zp & T==`Ttwo & phi1)
			 | (OP==`ADC_zp & T==`Ttwo & phi2)
			 | (OP==`ROR_zp & T==`Tzero & phi1)
			 | (OP==`ROR_zp & T==`Tzero & phi2)
			 | (OP==`ROR_zp & T==`Tone & phi1)
			 | (OP==`ROR_zp & T==`Tone & phi2)
			 | (OP==`ROR_zp & T==`Ttwo & phi1)
			 | (OP==`ROR_zp & T==`Ttwo & phi2)
			 | (OP==`ROR_zp & T==`Tthree & phi1)
			 | (OP==`ROR_zp & T==`Tthree & phi2)
			 | (OP==`ROR_zp & T==`Tfour & phi1)
			 | (OP==`ROR_zp & T==`Tfour & phi2)
			 | (OP==`PLA & T==`Tzero & phi1)
			 | (OP==`PLA & T==`Tzero & phi2)
			 | (OP==`PLA & T==`Tone & phi1)
			 | (OP==`PLA & T==`Tone & phi2)
			 | (OP==`PLA & T==`Ttwo & phi1)
			 | (OP==`PLA & T==`Ttwo & phi2)
			 | (OP==`PLA & T==`Tthree & phi1)
			 | (OP==`PLA & T==`Tthree & phi2)
			 | (OP==`ADC_imm & T==`Tone & phi1)
			 | (OP==`ADC_imm & T==`Tone & phi2)
			 | (OP==`ADC_imm & T==`Ttwo & phi1)
			 | (OP==`ADC_imm & T==`Ttwo & phi2)
			 | (OP==`ROR & T==`Tone & phi1)
			 | (OP==`ROR & T==`Tone & phi2)
			 | (OP==`ROR & T==`Ttwo & phi1)
			 | (OP==`ROR & T==`Ttwo & phi2)
			 | (OP==`JMP_zp & T==`Tzero & phi1)
			 | (OP==`JMP_zp & T==`Tzero & phi2)
			 | (OP==`JMP_zp & T==`Tone & phi1)
			 | (OP==`JMP_zp & T==`Tone & phi2)
			 | (OP==`JMP_zp & T==`Ttwo & phi1)
			 | (OP==`JMP_zp & T==`Ttwo & phi2)
			 | (OP==`JMP_zp & T==`Tthree & phi1)
			 | (OP==`JMP_zp & T==`Tthree & phi2)
			 | (OP==`JMP_zp & T==`Tfour & phi1)
			 | (OP==`JMP_zp & T==`Tfour & phi2)
			 | (OP==`ADC_abs & T==`Tzero & phi1)
			 | (OP==`ADC_abs & T==`Tzero & phi2)
			 | (OP==`ADC_abs & T==`Tone & phi1)
			 | (OP==`ADC_abs & T==`Tone & phi2)
			 | (OP==`ADC_abs & T==`Ttwo & phi1)
			 | (OP==`ADC_abs & T==`Ttwo & phi2)
			 | (OP==`ADC_abs & T==`Tthree & phi1)
			 | (OP==`ADC_abs & T==`Tthree & phi2)
			 | (OP==`ROR_abs & T==`Tzero & phi1)
			 | (OP==`ROR_abs & T==`Tzero & phi2)
			 | (OP==`ROR_abs & T==`Tone & phi1)
			 | (OP==`ROR_abs & T==`Tone & phi2)
			 | (OP==`ROR_abs & T==`Ttwo & phi1)
			 | (OP==`ROR_abs & T==`Ttwo & phi2)
			 | (OP==`ROR_abs & T==`Tthree & phi1)
			 | (OP==`ROR_abs & T==`Tthree & phi2)
			 | (OP==`ROR_abs & T==`Tfour & phi1)
			 | (OP==`ROR_abs & T==`Tfour & phi2)
			 | (OP==`ROR_abs & T==`Tfive & phi1)
			 | (OP==`ROR_abs & T==`Tfive & phi2)
			 | (OP==`BVS_rel & T==`Tzero & phi1)
			 | (OP==`BVS_rel & T==`Tzero & phi2)
			 | (OP==`BVS_rel & T==`Ttwo & phi1)
			 | (OP==`BVS_rel & T==`Ttwo & phi2)
			 | (OP==`BVS_rel & T==`Tthree & phi1)
			 | (OP==`BVS_rel & T==`Tthree & phi2)
			 | (OP==`BVS_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BVS_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BVS_rel & T==`T1BranchCross & phi1)
			 | (OP==`BVS_rel & T==`T1BranchCross & phi2)
			 | (OP==`BVS_rel & T==`T1NoBranch & phi1)
			 | (OP==`BVS_rel & T==`T1NoBranch & phi2)
			 | (OP==`ADC_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ADC_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`ADC_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`ADC_izy & T==`TzeroCrossPg & phi2)
			 | (OP==`ADC_izy & T==`Tone & phi1)
			 | (OP==`ADC_izy & T==`Tone & phi2)
			 | (OP==`ADC_izy & T==`Ttwo & phi1)
			 | (OP==`ADC_izy & T==`Ttwo & phi2)
			 | (OP==`ADC_izy & T==`Tthree & phi1)
			 | (OP==`ADC_izy & T==`Tthree & phi2)
			 | (OP==`ADC_izy & T==`Tfour & phi1)
			 | (OP==`ADC_izy & T==`Tfour & phi2)
			 | (OP==`ADC_izy & T==`Tfive & phi1)
			 | (OP==`ADC_izy & T==`Tfive & phi2)
			 | (OP==`ADC_zpx & T==`Tzero & phi1)
			 | (OP==`ADC_zpx & T==`Tzero & phi2)
			 | (OP==`ADC_zpx & T==`Tone & phi1)
			 | (OP==`ADC_zpx & T==`Tone & phi2)
			 | (OP==`ADC_zpx & T==`Ttwo & phi1)
			 | (OP==`ADC_zpx & T==`Ttwo & phi2)
			 | (OP==`ADC_zpx & T==`Tthree & phi1)
			 | (OP==`ADC_zpx & T==`Tthree & phi2)
			 | (OP==`ROR_zpx & T==`Tzero & phi1)
			 | (OP==`ROR_zpx & T==`Tzero & phi2)
			 | (OP==`ROR_zpx & T==`Tone & phi1)
			 | (OP==`ROR_zpx & T==`Tone & phi2)
			 | (OP==`ROR_zpx & T==`Ttwo & phi1)
			 | (OP==`ROR_zpx & T==`Ttwo & phi2)
			 | (OP==`ROR_zpx & T==`Tthree & phi1)
			 | (OP==`ROR_zpx & T==`Tthree & phi2)
			 | (OP==`ROR_zpx & T==`Tfour & phi1)
			 | (OP==`ROR_zpx & T==`Tfour & phi2)
			 | (OP==`ROR_zpx & T==`Tfive & phi1)
			 | (OP==`ROR_zpx & T==`Tfive & phi2)
			 | (OP==`SEI & T==`Tone & phi1)
			 | (OP==`SEI & T==`Tone & phi2)
			 | (OP==`SEI & T==`Ttwo & phi1)
			 | (OP==`SEI & T==`Ttwo & phi2)
			 | (OP==`ADC_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ADC_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`ADC_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`ADC_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`ADC_aby & T==`Tone & phi1)
			 | (OP==`ADC_aby & T==`Tone & phi2)
			 | (OP==`ADC_aby & T==`Ttwo & phi1)
			 | (OP==`ADC_aby & T==`Ttwo & phi2)
			 | (OP==`ADC_aby & T==`Tthree & phi1)
			 | (OP==`ADC_aby & T==`Tthree & phi2)
			 | (OP==`ADC_aby & T==`Tfour & phi1)
			 | (OP==`ADC_aby & T==`Tfour & phi2)
			 | (OP==`ADC_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ADC_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`ADC_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`ADC_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`ADC_abx & T==`Tone & phi1)
			 | (OP==`ADC_abx & T==`Tone & phi2)
			 | (OP==`ADC_abx & T==`Ttwo & phi1)
			 | (OP==`ADC_abx & T==`Ttwo & phi2)
			 | (OP==`ADC_abx & T==`Tthree & phi1)
			 | (OP==`ADC_abx & T==`Tthree & phi2)
			 | (OP==`ADC_abx & T==`Tfour & phi1)
			 | (OP==`ADC_abx & T==`Tfour & phi2)
			 | (OP==`ROR_abx & T==`Tzero & phi1)
			 | (OP==`ROR_abx & T==`Tzero & phi2)
			 | (OP==`ROR_abx & T==`Tone & phi1)
			 | (OP==`ROR_abx & T==`Tone & phi2)
			 | (OP==`ROR_abx & T==`Ttwo & phi1)
			 | (OP==`ROR_abx & T==`Ttwo & phi2)
			 | (OP==`ROR_abx & T==`Tthree & phi1)
			 | (OP==`ROR_abx & T==`Tthree & phi2)
			 | (OP==`ROR_abx & T==`Tfour & phi1)
			 | (OP==`ROR_abx & T==`Tfour & phi2)
			 | (OP==`ROR_abx & T==`Tfive & phi1)
			 | (OP==`ROR_abx & T==`Tfive & phi2)
			 | (OP==`ROR_abx & T==`Tsix & phi1)
			 | (OP==`ROR_abx & T==`Tsix & phi2)
			 | (OP==`STA_izx & T==`Tzero & phi1)
			 | (OP==`STA_izx & T==`Tzero & phi2)
			 | (OP==`STA_izx & T==`Tone & phi1)
			 | (OP==`STA_izx & T==`Tone & phi2)
			 | (OP==`STA_izx & T==`Ttwo & phi1)
			 | (OP==`STA_izx & T==`Ttwo & phi2)
			 | (OP==`STA_izx & T==`Tthree & phi1)
			 | (OP==`STA_izx & T==`Tthree & phi2)
			 | (OP==`STA_izx & T==`Tfour & phi1)
			 | (OP==`STA_izx & T==`Tfour & phi2)
			 | (OP==`STA_izx & T==`Tfive & phi1)
			 | (OP==`STA_izx & T==`Tfive & phi2)
			 | (OP==`STY_zp & T==`Tzero & phi1)
			 | (OP==`STY_zp & T==`Tzero & phi2)
			 | (OP==`STY_zp & T==`Tone & phi1)
			 | (OP==`STY_zp & T==`Tone & phi2)
			 | (OP==`STY_zp & T==`Ttwo & phi1)
			 | (OP==`STY_zp & T==`Ttwo & phi2)
			 | (OP==`STA_zp & T==`Tzero & phi1)
			 | (OP==`STA_zp & T==`Tzero & phi2)
			 | (OP==`STA_zp & T==`Tone & phi1)
			 | (OP==`STA_zp & T==`Tone & phi2)
			 | (OP==`STA_zp & T==`Ttwo & phi1)
			 | (OP==`STA_zp & T==`Ttwo & phi2)
			 | (OP==`STX_zp & T==`Tzero & phi1)
			 | (OP==`STX_zp & T==`Tzero & phi2)
			 | (OP==`STX_zp & T==`Tone & phi1)
			 | (OP==`STX_zp & T==`Tone & phi2)
			 | (OP==`STX_zp & T==`Ttwo & phi1)
			 | (OP==`STX_zp & T==`Ttwo & phi2)
			 | (OP==`DEY & T==`Tone & phi1)
			 | (OP==`DEY & T==`Tone & phi2)
			 | (OP==`DEY & T==`Ttwo & phi1)
			 | (OP==`DEY & T==`Ttwo & phi2)
			 | (OP==`TXA & T==`Tone & phi1)
			 | (OP==`TXA & T==`Tone & phi2)
			 | (OP==`TXA & T==`Ttwo & phi1)
			 | (OP==`TXA & T==`Ttwo & phi2)
			 | (OP==`STY_abs & T==`Tzero & phi1)
			 | (OP==`STY_abs & T==`Tzero & phi2)
			 | (OP==`STY_abs & T==`Tone & phi1)
			 | (OP==`STY_abs & T==`Tone & phi2)
			 | (OP==`STY_abs & T==`Ttwo & phi1)
			 | (OP==`STY_abs & T==`Ttwo & phi2)
			 | (OP==`STY_abs & T==`Tthree & phi1)
			 | (OP==`STY_abs & T==`Tthree & phi2)
			 | (OP==`STA_abs & T==`Tzero & phi1)
			 | (OP==`STA_abs & T==`Tzero & phi2)
			 | (OP==`STA_abs & T==`Tone & phi1)
			 | (OP==`STA_abs & T==`Tone & phi2)
			 | (OP==`STA_abs & T==`Ttwo & phi1)
			 | (OP==`STA_abs & T==`Ttwo & phi2)
			 | (OP==`STA_abs & T==`Tthree & phi1)
			 | (OP==`STA_abs & T==`Tthree & phi2)
			 | (OP==`STX_abs & T==`Tzero & phi1)
			 | (OP==`STX_abs & T==`Tzero & phi2)
			 | (OP==`STX_abs & T==`Tone & phi1)
			 | (OP==`STX_abs & T==`Tone & phi2)
			 | (OP==`STX_abs & T==`Ttwo & phi1)
			 | (OP==`STX_abs & T==`Ttwo & phi2)
			 | (OP==`STX_abs & T==`Tthree & phi1)
			 | (OP==`STX_abs & T==`Tthree & phi2)
			 | (OP==`BCC_rel & T==`Tzero & phi1)
			 | (OP==`BCC_rel & T==`Tzero & phi2)
			 | (OP==`BCC_rel & T==`Ttwo & phi1)
			 | (OP==`BCC_rel & T==`Ttwo & phi2)
			 | (OP==`BCC_rel & T==`Tthree & phi1)
			 | (OP==`BCC_rel & T==`Tthree & phi2)
			 | (OP==`BCC_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BCC_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BCC_rel & T==`T1BranchCross & phi1)
			 | (OP==`BCC_rel & T==`T1BranchCross & phi2)
			 | (OP==`BCC_rel & T==`T1NoBranch & phi1)
			 | (OP==`BCC_rel & T==`T1NoBranch & phi2)
			 | (OP==`STA_izy & T==`Tzero & phi1)
			 | (OP==`STA_izy & T==`Tzero & phi2)
			 | (OP==`STA_izy & T==`Tone & phi1)
			 | (OP==`STA_izy & T==`Tone & phi2)
			 | (OP==`STA_izy & T==`Ttwo & phi1)
			 | (OP==`STA_izy & T==`Ttwo & phi2)
			 | (OP==`STA_izy & T==`Tthree & phi1)
			 | (OP==`STA_izy & T==`Tthree & phi2)
			 | (OP==`STA_izy & T==`Tfour & phi1)
			 | (OP==`STA_izy & T==`Tfour & phi2)
			 | (OP==`STA_izy & T==`Tfive & phi1)
			 | (OP==`STA_izy & T==`Tfive & phi2)
			 | (OP==`STY_zpx & T==`Tzero & phi1)
			 | (OP==`STY_zpx & T==`Tzero & phi2)
			 | (OP==`STY_zpx & T==`Tone & phi1)
			 | (OP==`STY_zpx & T==`Tone & phi2)
			 | (OP==`STY_zpx & T==`Ttwo & phi1)
			 | (OP==`STY_zpx & T==`Ttwo & phi2)
			 | (OP==`STY_zpx & T==`Tthree & phi1)
			 | (OP==`STY_zpx & T==`Tthree & phi2)
			 | (OP==`STA_zpx & T==`Tzero & phi1)
			 | (OP==`STA_zpx & T==`Tzero & phi2)
			 | (OP==`STA_zpx & T==`Tone & phi1)
			 | (OP==`STA_zpx & T==`Tone & phi2)
			 | (OP==`STA_zpx & T==`Ttwo & phi1)
			 | (OP==`STA_zpx & T==`Ttwo & phi2)
			 | (OP==`STA_zpx & T==`Tthree & phi1)
			 | (OP==`STA_zpx & T==`Tthree & phi2)
			 | (OP==`STX_zpy & T==`Tzero & phi1)
			 | (OP==`STX_zpy & T==`Tzero & phi2)
			 | (OP==`STX_zpy & T==`Tone & phi1)
			 | (OP==`STX_zpy & T==`Tone & phi2)
			 | (OP==`STX_zpy & T==`Ttwo & phi1)
			 | (OP==`STX_zpy & T==`Ttwo & phi2)
			 | (OP==`STX_zpy & T==`Tthree & phi1)
			 | (OP==`STX_zpy & T==`Tthree & phi2)
			 | (OP==`TYA & T==`Tone & phi1)
			 | (OP==`TYA & T==`Tone & phi2)
			 | (OP==`TYA & T==`Ttwo & phi1)
			 | (OP==`TYA & T==`Ttwo & phi2)
			 | (OP==`STA_aby & T==`Tzero & phi1)
			 | (OP==`STA_aby & T==`Tzero & phi2)
			 | (OP==`STA_aby & T==`Tone & phi1)
			 | (OP==`STA_aby & T==`Tone & phi2)
			 | (OP==`STA_aby & T==`Ttwo & phi1)
			 | (OP==`STA_aby & T==`Ttwo & phi2)
			 | (OP==`STA_aby & T==`Tthree & phi1)
			 | (OP==`STA_aby & T==`Tthree & phi2)
			 | (OP==`STA_aby & T==`Tfour & phi1)
			 | (OP==`STA_aby & T==`Tfour & phi2)
			 | (OP==`TXS & T==`Tone & phi1)
			 | (OP==`TXS & T==`Tone & phi2)
			 | (OP==`TXS & T==`Ttwo & phi1)
			 | (OP==`TXS & T==`Ttwo & phi2)
			 | (OP==`STA_abx & T==`Tzero & phi1)
			 | (OP==`STA_abx & T==`Tzero & phi2)
			 | (OP==`STA_abx & T==`Tone & phi1)
			 | (OP==`STA_abx & T==`Tone & phi2)
			 | (OP==`STA_abx & T==`Ttwo & phi1)
			 | (OP==`STA_abx & T==`Ttwo & phi2)
			 | (OP==`STA_abx & T==`Tthree & phi1)
			 | (OP==`STA_abx & T==`Tthree & phi2)
			 | (OP==`STA_abx & T==`Tfour & phi1)
			 | (OP==`STA_abx & T==`Tfour & phi2)
			 | (OP==`LDY_imm & T==`Tone & phi1)
			 | (OP==`LDY_imm & T==`Tone & phi2)
			 | (OP==`LDY_imm & T==`Ttwo & phi1)
			 | (OP==`LDY_imm & T==`Ttwo & phi2)
			 | (OP==`LDA_izx & T==`Tzero & phi1)
			 | (OP==`LDA_izx & T==`Tzero & phi2)
			 | (OP==`LDA_izx & T==`Tone & phi1)
			 | (OP==`LDA_izx & T==`Tone & phi2)
			 | (OP==`LDA_izx & T==`Ttwo & phi1)
			 | (OP==`LDA_izx & T==`Ttwo & phi2)
			 | (OP==`LDA_izx & T==`Tthree & phi1)
			 | (OP==`LDA_izx & T==`Tthree & phi2)
			 | (OP==`LDA_izx & T==`Tfour & phi1)
			 | (OP==`LDA_izx & T==`Tfour & phi2)
			 | (OP==`LDA_izx & T==`Tfive & phi1)
			 | (OP==`LDA_izx & T==`Tfive & phi2)
			 | (OP==`LDX_imm & T==`Tone & phi1)
			 | (OP==`LDX_imm & T==`Tone & phi2)
			 | (OP==`LDX_imm & T==`Ttwo & phi1)
			 | (OP==`LDX_imm & T==`Ttwo & phi2)
			 | (OP==`LDY_zp & T==`Tzero & phi1)
			 | (OP==`LDY_zp & T==`Tzero & phi2)
			 | (OP==`LDY_zp & T==`Tone & phi1)
			 | (OP==`LDY_zp & T==`Tone & phi2)
			 | (OP==`LDY_zp & T==`Ttwo & phi1)
			 | (OP==`LDY_zp & T==`Ttwo & phi2)
			 | (OP==`LDA_zp & T==`Tzero & phi1)
			 | (OP==`LDA_zp & T==`Tzero & phi2)
			 | (OP==`LDA_zp & T==`Tone & phi1)
			 | (OP==`LDA_zp & T==`Tone & phi2)
			 | (OP==`LDA_zp & T==`Ttwo & phi1)
			 | (OP==`LDA_zp & T==`Ttwo & phi2)
			 | (OP==`LDX_zp & T==`Tzero & phi1)
			 | (OP==`LDX_zp & T==`Tzero & phi2)
			 | (OP==`LDX_zp & T==`Tone & phi1)
			 | (OP==`LDX_zp & T==`Tone & phi2)
			 | (OP==`LDX_zp & T==`Ttwo & phi1)
			 | (OP==`LDX_zp & T==`Ttwo & phi2)
			 | (OP==`TAY & T==`Tone & phi1)
			 | (OP==`TAY & T==`Tone & phi2)
			 | (OP==`TAY & T==`Ttwo & phi1)
			 | (OP==`TAY & T==`Ttwo & phi2)
			 | (OP==`LDA_imm & T==`Tone & phi1)
			 | (OP==`LDA_imm & T==`Tone & phi2)
			 | (OP==`LDA_imm & T==`Ttwo & phi1)
			 | (OP==`LDA_imm & T==`Ttwo & phi2)
			 | (OP==`TAX & T==`Tone & phi1)
			 | (OP==`TAX & T==`Tone & phi2)
			 | (OP==`TAX & T==`Ttwo & phi1)
			 | (OP==`TAX & T==`Ttwo & phi2)
			 | (OP==`LDY_abs & T==`Tzero & phi1)
			 | (OP==`LDY_abs & T==`Tzero & phi2)
			 | (OP==`LDY_abs & T==`Tone & phi1)
			 | (OP==`LDY_abs & T==`Tone & phi2)
			 | (OP==`LDY_abs & T==`Ttwo & phi1)
			 | (OP==`LDY_abs & T==`Ttwo & phi2)
			 | (OP==`LDY_abs & T==`Tthree & phi1)
			 | (OP==`LDY_abs & T==`Tthree & phi2)
			 | (OP==`LDA_abs & T==`Tzero & phi1)
			 | (OP==`LDA_abs & T==`Tzero & phi2)
			 | (OP==`LDA_abs & T==`Tone & phi1)
			 | (OP==`LDA_abs & T==`Tone & phi2)
			 | (OP==`LDA_abs & T==`Ttwo & phi1)
			 | (OP==`LDA_abs & T==`Ttwo & phi2)
			 | (OP==`LDA_abs & T==`Tthree & phi1)
			 | (OP==`LDA_abs & T==`Tthree & phi2)
			 | (OP==`LDX_abs & T==`Tzero & phi1)
			 | (OP==`LDX_abs & T==`Tzero & phi2)
			 | (OP==`LDX_abs & T==`Tone & phi1)
			 | (OP==`LDX_abs & T==`Tone & phi2)
			 | (OP==`LDX_abs & T==`Ttwo & phi1)
			 | (OP==`LDX_abs & T==`Ttwo & phi2)
			 | (OP==`LDX_abs & T==`Tthree & phi1)
			 | (OP==`LDX_abs & T==`Tthree & phi2)
			 | (OP==`BCS_rel & T==`Tzero & phi1)
			 | (OP==`BCS_rel & T==`Tzero & phi2)
			 | (OP==`BCS_rel & T==`Ttwo & phi1)
			 | (OP==`BCS_rel & T==`Ttwo & phi2)
			 | (OP==`BCS_rel & T==`Tthree & phi1)
			 | (OP==`BCS_rel & T==`Tthree & phi2)
			 | (OP==`BCS_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BCS_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BCS_rel & T==`T1BranchCross & phi1)
			 | (OP==`BCS_rel & T==`T1BranchCross & phi2)
			 | (OP==`BCS_rel & T==`T1NoBranch & phi1)
			 | (OP==`BCS_rel & T==`T1NoBranch & phi2)
			 | (OP==`LDA_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDA_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`LDA_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`LDA_izy & T==`TzeroCrossPg & phi2)
			 | (OP==`LDA_izy & T==`Tone & phi1)
			 | (OP==`LDA_izy & T==`Tone & phi2)
			 | (OP==`LDA_izy & T==`Ttwo & phi1)
			 | (OP==`LDA_izy & T==`Ttwo & phi2)
			 | (OP==`LDA_izy & T==`Tthree & phi1)
			 | (OP==`LDA_izy & T==`Tthree & phi2)
			 | (OP==`LDA_izy & T==`Tfour & phi1)
			 | (OP==`LDA_izy & T==`Tfour & phi2)
			 | (OP==`LDA_izy & T==`Tfive & phi1)
			 | (OP==`LDA_izy & T==`Tfive & phi2)
			 | (OP==`LDY_zpx & T==`Tzero & phi1)
			 | (OP==`LDY_zpx & T==`Tzero & phi2)
			 | (OP==`LDY_zpx & T==`Tone & phi1)
			 | (OP==`LDY_zpx & T==`Tone & phi2)
			 | (OP==`LDY_zpx & T==`Ttwo & phi1)
			 | (OP==`LDY_zpx & T==`Ttwo & phi2)
			 | (OP==`LDY_zpx & T==`Tthree & phi1)
			 | (OP==`LDY_zpx & T==`Tthree & phi2)
			 | (OP==`LDA_zpx & T==`Tzero & phi1)
			 | (OP==`LDA_zpx & T==`Tzero & phi2)
			 | (OP==`LDA_zpx & T==`Tone & phi1)
			 | (OP==`LDA_zpx & T==`Tone & phi2)
			 | (OP==`LDA_zpx & T==`Ttwo & phi1)
			 | (OP==`LDA_zpx & T==`Ttwo & phi2)
			 | (OP==`LDA_zpx & T==`Tthree & phi1)
			 | (OP==`LDA_zpx & T==`Tthree & phi2)
			 | (OP==`LDX_zpy & T==`Tzero & phi1)
			 | (OP==`LDX_zpy & T==`Tzero & phi2)
			 | (OP==`LDX_zpy & T==`Tone & phi1)
			 | (OP==`LDX_zpy & T==`Tone & phi2)
			 | (OP==`LDX_zpy & T==`Ttwo & phi1)
			 | (OP==`LDX_zpy & T==`Ttwo & phi2)
			 | (OP==`LDX_zpy & T==`Tthree & phi1)
			 | (OP==`LDX_zpy & T==`Tthree & phi2)
			 | (OP==`CLV & T==`Tone & phi1)
			 | (OP==`CLV & T==`Tone & phi2)
			 | (OP==`CLV & T==`Ttwo & phi1)
			 | (OP==`CLV & T==`Ttwo & phi2)
			 | (OP==`LDA_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDA_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`LDA_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`LDA_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`LDA_aby & T==`Tone & phi1)
			 | (OP==`LDA_aby & T==`Tone & phi2)
			 | (OP==`LDA_aby & T==`Ttwo & phi1)
			 | (OP==`LDA_aby & T==`Ttwo & phi2)
			 | (OP==`LDA_aby & T==`Tthree & phi1)
			 | (OP==`LDA_aby & T==`Tthree & phi2)
			 | (OP==`LDA_aby & T==`Tfour & phi1)
			 | (OP==`LDA_aby & T==`Tfour & phi2)
			 | (OP==`TSX & T==`Tone & phi1)
			 | (OP==`TSX & T==`Tone & phi2)
			 | (OP==`TSX & T==`Ttwo & phi1)
			 | (OP==`TSX & T==`Ttwo & phi2)
			 | (OP==`LDY_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDY_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`LDY_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`LDY_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`LDY_abx & T==`Tone & phi1)
			 | (OP==`LDY_abx & T==`Tone & phi2)
			 | (OP==`LDY_abx & T==`Ttwo & phi1)
			 | (OP==`LDY_abx & T==`Ttwo & phi2)
			 | (OP==`LDY_abx & T==`Tthree & phi1)
			 | (OP==`LDY_abx & T==`Tthree & phi2)
			 | (OP==`LDY_abx & T==`Tfour & phi1)
			 | (OP==`LDY_abx & T==`Tfour & phi2)
			 | (OP==`LDA_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDA_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`LDA_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`LDA_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`LDA_abx & T==`Tone & phi1)
			 | (OP==`LDA_abx & T==`Tone & phi2)
			 | (OP==`LDA_abx & T==`Ttwo & phi1)
			 | (OP==`LDA_abx & T==`Ttwo & phi2)
			 | (OP==`LDA_abx & T==`Tthree & phi1)
			 | (OP==`LDA_abx & T==`Tthree & phi2)
			 | (OP==`LDA_abx & T==`Tfour & phi1)
			 | (OP==`LDA_abx & T==`Tfour & phi2)
			 | (OP==`LDX_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDX_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`LDX_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`LDX_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`LDX_aby & T==`Tone & phi1)
			 | (OP==`LDX_aby & T==`Tone & phi2)
			 | (OP==`LDX_aby & T==`Ttwo & phi1)
			 | (OP==`LDX_aby & T==`Ttwo & phi2)
			 | (OP==`LDX_aby & T==`Tthree & phi1)
			 | (OP==`LDX_aby & T==`Tthree & phi2)
			 | (OP==`LDX_aby & T==`Tfour & phi1)
			 | (OP==`LDX_aby & T==`Tfour & phi2)
			 | (OP==`CPY_imm & T==`Tone & phi1)
			 | (OP==`CPY_imm & T==`Tone & phi2)
			 | (OP==`CPY_imm & T==`Ttwo & phi1)
			 | (OP==`CPY_imm & T==`Ttwo & phi2)
			 | (OP==`CMP_izx & T==`Tzero & phi1)
			 | (OP==`CMP_izx & T==`Tzero & phi2)
			 | (OP==`CMP_izx & T==`Tone & phi1)
			 | (OP==`CMP_izx & T==`Tone & phi2)
			 | (OP==`CMP_izx & T==`Ttwo & phi1)
			 | (OP==`CMP_izx & T==`Ttwo & phi2)
			 | (OP==`CMP_izx & T==`Tthree & phi1)
			 | (OP==`CMP_izx & T==`Tthree & phi2)
			 | (OP==`CMP_izx & T==`Tfour & phi1)
			 | (OP==`CMP_izx & T==`Tfour & phi2)
			 | (OP==`CMP_izx & T==`Tfive & phi1)
			 | (OP==`CMP_izx & T==`Tfive & phi2)
			 | (OP==`CPY_zp & T==`Tzero & phi1)
			 | (OP==`CPY_zp & T==`Tzero & phi2)
			 | (OP==`CPY_zp & T==`Tone & phi1)
			 | (OP==`CPY_zp & T==`Tone & phi2)
			 | (OP==`CPY_zp & T==`Ttwo & phi1)
			 | (OP==`CPY_zp & T==`Ttwo & phi2)
			 | (OP==`CMP_zp & T==`Tzero & phi1)
			 | (OP==`CMP_zp & T==`Tzero & phi2)
			 | (OP==`CMP_zp & T==`Tone & phi1)
			 | (OP==`CMP_zp & T==`Tone & phi2)
			 | (OP==`CMP_zp & T==`Ttwo & phi1)
			 | (OP==`CMP_zp & T==`Ttwo & phi2)
			 | (OP==`DEC_zp & T==`Tzero & phi1)
			 | (OP==`DEC_zp & T==`Tzero & phi2)
			 | (OP==`DEC_zp & T==`Tone & phi1)
			 | (OP==`DEC_zp & T==`Tone & phi2)
			 | (OP==`DEC_zp & T==`Ttwo & phi1)
			 | (OP==`DEC_zp & T==`Ttwo & phi2)
			 | (OP==`DEC_zp & T==`Tthree & phi1)
			 | (OP==`DEC_zp & T==`Tthree & phi2)
			 | (OP==`DEC_zp & T==`Tfour & phi1)
			 | (OP==`DEC_zp & T==`Tfour & phi2)
			 | (OP==`INY & T==`Tone & phi1)
			 | (OP==`INY & T==`Tone & phi2)
			 | (OP==`INY & T==`Ttwo & phi1)
			 | (OP==`INY & T==`Ttwo & phi2)
			 | (OP==`CMP_imm & T==`Tone & phi1)
			 | (OP==`CMP_imm & T==`Tone & phi2)
			 | (OP==`CMP_imm & T==`Ttwo & phi1)
			 | (OP==`CMP_imm & T==`Ttwo & phi2)
			 | (OP==`DEX & T==`Tone & phi1)
			 | (OP==`DEX & T==`Tone & phi2)
			 | (OP==`DEX & T==`Ttwo & phi1)
			 | (OP==`DEX & T==`Ttwo & phi2)
			 | (OP==`CPY_abs & T==`Tzero & phi1)
			 | (OP==`CPY_abs & T==`Tzero & phi2)
			 | (OP==`CPY_abs & T==`Tone & phi1)
			 | (OP==`CPY_abs & T==`Tone & phi2)
			 | (OP==`CPY_abs & T==`Ttwo & phi1)
			 | (OP==`CPY_abs & T==`Ttwo & phi2)
			 | (OP==`CPY_abs & T==`Tthree & phi1)
			 | (OP==`CPY_abs & T==`Tthree & phi2)
			 | (OP==`CMP_abs & T==`Tzero & phi1)
			 | (OP==`CMP_abs & T==`Tzero & phi2)
			 | (OP==`CMP_abs & T==`Tone & phi1)
			 | (OP==`CMP_abs & T==`Tone & phi2)
			 | (OP==`CMP_abs & T==`Ttwo & phi1)
			 | (OP==`CMP_abs & T==`Ttwo & phi2)
			 | (OP==`CMP_abs & T==`Tthree & phi1)
			 | (OP==`CMP_abs & T==`Tthree & phi2)
			 | (OP==`DEC_abs & T==`Tzero & phi1)
			 | (OP==`DEC_abs & T==`Tzero & phi2)
			 | (OP==`DEC_abs & T==`Tone & phi1)
			 | (OP==`DEC_abs & T==`Tone & phi2)
			 | (OP==`DEC_abs & T==`Ttwo & phi1)
			 | (OP==`DEC_abs & T==`Ttwo & phi2)
			 | (OP==`DEC_abs & T==`Tthree & phi1)
			 | (OP==`DEC_abs & T==`Tthree & phi2)
			 | (OP==`DEC_abs & T==`Tfour & phi1)
			 | (OP==`DEC_abs & T==`Tfour & phi2)
			 | (OP==`DEC_abs & T==`Tfive & phi1)
			 | (OP==`DEC_abs & T==`Tfive & phi2)
			 | (OP==`BNE_rel & T==`Tzero & phi1)
			 | (OP==`BNE_rel & T==`Tzero & phi2)
			 | (OP==`BNE_rel & T==`Ttwo & phi1)
			 | (OP==`BNE_rel & T==`Ttwo & phi2)
			 | (OP==`BNE_rel & T==`Tthree & phi1)
			 | (OP==`BNE_rel & T==`Tthree & phi2)
			 | (OP==`BNE_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BNE_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BNE_rel & T==`T1BranchCross & phi1)
			 | (OP==`BNE_rel & T==`T1BranchCross & phi2)
			 | (OP==`BNE_rel & T==`T1NoBranch & phi1)
			 | (OP==`BNE_rel & T==`T1NoBranch & phi2)
			 | (OP==`CMP_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`CMP_izy & T==`TzeroCrossPg & phi2)
			 | (OP==`CMP_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`CMP_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`CMP_izy & T==`Tone & phi1)
			 | (OP==`CMP_izy & T==`Tone & phi2)
			 | (OP==`CMP_izy & T==`Ttwo & phi1)
			 | (OP==`CMP_izy & T==`Ttwo & phi2)
			 | (OP==`CMP_izy & T==`Tthree & phi1)
			 | (OP==`CMP_izy & T==`Tthree & phi2)
			 | (OP==`CMP_izy & T==`Tfour & phi1)
			 | (OP==`CMP_izy & T==`Tfour & phi2)
			 | (OP==`CMP_izy & T==`Tfive & phi1)
			 | (OP==`CMP_izy & T==`Tfive & phi2)
			 | (OP==`CMP_zpx & T==`Tzero & phi1)
			 | (OP==`CMP_zpx & T==`Tzero & phi2)
			 | (OP==`CMP_zpx & T==`Tone & phi1)
			 | (OP==`CMP_zpx & T==`Tone & phi2)
			 | (OP==`CMP_zpx & T==`Ttwo & phi1)
			 | (OP==`CMP_zpx & T==`Ttwo & phi2)
			 | (OP==`CMP_zpx & T==`Tthree & phi1)
			 | (OP==`CMP_zpx & T==`Tthree & phi2)
			 | (OP==`DEC_zpx & T==`Tzero & phi1)
			 | (OP==`DEC_zpx & T==`Tzero & phi2)
			 | (OP==`DEC_zpx & T==`Tone & phi1)
			 | (OP==`DEC_zpx & T==`Tone & phi2)
			 | (OP==`DEC_zpx & T==`Ttwo & phi1)
			 | (OP==`DEC_zpx & T==`Ttwo & phi2)
			 | (OP==`DEC_zpx & T==`Tthree & phi1)
			 | (OP==`DEC_zpx & T==`Tthree & phi2)
			 | (OP==`DEC_zpx & T==`Tfour & phi1)
			 | (OP==`DEC_zpx & T==`Tfour & phi2)
			 | (OP==`DEC_zpx & T==`Tfive & phi1)
			 | (OP==`DEC_zpx & T==`Tfive & phi2)
			 | (OP==`CLD & T==`Tone & phi1)
			 | (OP==`CLD & T==`Tone & phi2)
			 | (OP==`CLD & T==`Ttwo & phi1)
			 | (OP==`CLD & T==`Ttwo & phi2)
			 | (OP==`CMP_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`CMP_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`CMP_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`CMP_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`CMP_aby & T==`Tone & phi1)
			 | (OP==`CMP_aby & T==`Tone & phi2)
			 | (OP==`CMP_aby & T==`Ttwo & phi1)
			 | (OP==`CMP_aby & T==`Ttwo & phi2)
			 | (OP==`CMP_aby & T==`Tthree & phi1)
			 | (OP==`CMP_aby & T==`Tthree & phi2)
			 | (OP==`CMP_aby & T==`Tfour & phi1)
			 | (OP==`CMP_aby & T==`Tfour & phi2)
			 | (OP==`CMP_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`CMP_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`CMP_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`CMP_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`CMP_abx & T==`Tone & phi1)
			 | (OP==`CMP_abx & T==`Tone & phi2)
			 | (OP==`CMP_abx & T==`Ttwo & phi1)
			 | (OP==`CMP_abx & T==`Ttwo & phi2)
			 | (OP==`CMP_abx & T==`Tthree & phi1)
			 | (OP==`CMP_abx & T==`Tthree & phi2)
			 | (OP==`CMP_abx & T==`Tfour & phi1)
			 | (OP==`CMP_abx & T==`Tfour & phi2)
			 | (OP==`DEC_abx & T==`Tzero & phi1)
			 | (OP==`DEC_abx & T==`Tzero & phi2)
			 | (OP==`DEC_abx & T==`Tone & phi1)
			 | (OP==`DEC_abx & T==`Tone & phi2)
			 | (OP==`DEC_abx & T==`Ttwo & phi1)
			 | (OP==`DEC_abx & T==`Ttwo & phi2)
			 | (OP==`DEC_abx & T==`Tthree & phi1)
			 | (OP==`DEC_abx & T==`Tthree & phi2)
			 | (OP==`DEC_abx & T==`Tfour & phi1)
			 | (OP==`DEC_abx & T==`Tfour & phi2)
			 | (OP==`DEC_abx & T==`Tfive & phi1)
			 | (OP==`DEC_abx & T==`Tfive & phi2)
			 | (OP==`DEC_abx & T==`Tsix & phi1)
			 | (OP==`DEC_abx & T==`Tsix & phi2)
			 | (OP==`CPX_imm & T==`Tone & phi1)
			 | (OP==`CPX_imm & T==`Tone & phi2)
			 | (OP==`CPX_imm & T==`Ttwo & phi1)
			 | (OP==`CPX_imm & T==`Ttwo & phi2)
			 | (OP==`SBC_izx & T==`Tzero & phi1)
			 | (OP==`SBC_izx & T==`Tzero & phi2)
			 | (OP==`SBC_izx & T==`Tone & phi1 & !decMode)
			 | (OP==`SBC_izx & T==`Tone & phi2 & !decMode)
			 | (OP==`SBC_izx & T==`Ttwo & phi1)
			 | (OP==`SBC_izx & T==`Ttwo & phi2)
			 | (OP==`SBC_izx & T==`Tthree & phi1)
			 | (OP==`SBC_izx & T==`Tthree & phi2)
			 | (OP==`SBC_izx & T==`Tfour & phi1)
			 | (OP==`SBC_izx & T==`Tfour & phi2)
			 | (OP==`SBC_izx & T==`Tfive & phi1)
			 | (OP==`SBC_izx & T==`Tfive & phi2)
			 | (OP==`CPX_zp & T==`Tzero & phi1)
			 | (OP==`CPX_zp & T==`Tzero & phi2)
			 | (OP==`CPX_zp & T==`Tone & phi1)
			 | (OP==`CPX_zp & T==`Tone & phi2)
			 | (OP==`CPX_zp & T==`Ttwo & phi1)
			 | (OP==`CPX_zp & T==`Ttwo & phi2)
			 | (OP==`SBC_zp & T==`Tzero & phi1)
			 | (OP==`SBC_zp & T==`Tzero & phi2)
			 | (OP==`SBC_zp & T==`Tone & phi1 & !decMode)
			 | (OP==`SBC_zp & T==`Tone & phi2 & !decMode)
			 | (OP==`SBC_zp & T==`Ttwo & phi1)
			 | (OP==`SBC_zp & T==`Ttwo & phi2)
			 | (OP==`INC_zp & T==`Tzero & phi1)
			 | (OP==`INC_zp & T==`Tzero & phi2)
			 | (OP==`INC_zp & T==`Tone & phi1)
			 | (OP==`INC_zp & T==`Tone & phi2)
			 | (OP==`INC_zp & T==`Ttwo & phi1)
			 | (OP==`INC_zp & T==`Ttwo & phi2)
			 | (OP==`INC_zp & T==`Tthree & phi1)
			 | (OP==`INC_zp & T==`Tthree & phi2)
			 | (OP==`INC_zp & T==`Tfour & phi1)
			 | (OP==`INC_zp & T==`Tfour & phi2)
			 | (OP==`INX & T==`Tone & phi1)
			 | (OP==`INX & T==`Tone & phi2)
			 | (OP==`INX & T==`Ttwo & phi1)
			 | (OP==`INX & T==`Ttwo & phi2)
			 | (OP==`SBC_imm & T==`Tone & phi1 & !decMode)
			 | (OP==`SBC_imm & T==`Tone & phi2 & !decMode)
			 | (OP==`SBC_imm & T==`Ttwo & phi1)
			 | (OP==`SBC_imm & T==`Ttwo & phi2)
			 | (OP==`NOP & T==`Tone & phi1)
			 | (OP==`NOP & T==`Tone & phi2)
			 | (OP==`NOP & T==`Ttwo & phi1)
			 | (OP==`NOP & T==`Ttwo & phi2)
			 | (OP==`CPX_abs & T==`Tzero & phi1)
			 | (OP==`CPX_abs & T==`Tzero & phi2)
			 | (OP==`CPX_abs & T==`Tone & phi1)
			 | (OP==`CPX_abs & T==`Tone & phi2)
			 | (OP==`CPX_abs & T==`Ttwo & phi1)
			 | (OP==`CPX_abs & T==`Ttwo & phi2)
			 | (OP==`CPX_abs & T==`Tthree & phi1)
			 | (OP==`CPX_abs & T==`Tthree & phi2)
			 | (OP==`SBC_abs & T==`Tzero & phi1)
			 | (OP==`SBC_abs & T==`Tzero & phi2)
			 | (OP==`SBC_abs & T==`Tone & phi1 & !decMode)
			 | (OP==`SBC_abs & T==`Tone & phi2 & !decMode)
			 | (OP==`SBC_abs & T==`Ttwo & phi1)
			 | (OP==`SBC_abs & T==`Ttwo & phi2)
			 | (OP==`SBC_abs & T==`Tthree & phi1)
			 | (OP==`SBC_abs & T==`Tthree & phi2)
			 | (OP==`INC_abs & T==`Tzero & phi1)
			 | (OP==`INC_abs & T==`Tzero & phi2)
			 | (OP==`INC_abs & T==`Tone & phi1)
			 | (OP==`INC_abs & T==`Tone & phi2)
			 | (OP==`INC_abs & T==`Ttwo & phi1)
			 | (OP==`INC_abs & T==`Ttwo & phi2)
			 | (OP==`INC_abs & T==`Tthree & phi1)
			 | (OP==`INC_abs & T==`Tthree & phi2)
			 | (OP==`INC_abs & T==`Tfour & phi1)
			 | (OP==`INC_abs & T==`Tfour & phi2)
			 | (OP==`INC_abs & T==`Tfive & phi1)
			 | (OP==`INC_abs & T==`Tfive & phi2)
			 | (OP==`BEQ_rel & T==`Tzero & phi1)
			 | (OP==`BEQ_rel & T==`Tzero & phi2)
			 | (OP==`BEQ_rel & T==`Ttwo & phi1)
			 | (OP==`BEQ_rel & T==`Ttwo & phi2)
			 | (OP==`BEQ_rel & T==`Tthree & phi1)
			 | (OP==`BEQ_rel & T==`Tthree & phi2)
			 | (OP==`BEQ_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BEQ_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BEQ_rel & T==`T1BranchCross & phi1)
			 | (OP==`BEQ_rel & T==`T1BranchCross & phi2)
			 | (OP==`BEQ_rel & T==`T1NoBranch & phi1)
			 | (OP==`BEQ_rel & T==`T1NoBranch & phi2)
			 | (OP==`SBC_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`SBC_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`SBC_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`SBC_izy & T==`TzeroCrossPg & phi2)
			 | (OP==`SBC_izy & T==`Tone & phi1 & !decMode)
			 | (OP==`SBC_izy & T==`Tone & phi2 & !decMode)
			 | (OP==`SBC_izy & T==`Ttwo & phi1)
			 | (OP==`SBC_izy & T==`Ttwo & phi2)
			 | (OP==`SBC_izy & T==`Tthree & phi1)
			 | (OP==`SBC_izy & T==`Tthree & phi2)
			 | (OP==`SBC_izy & T==`Tfour & phi1)
			 | (OP==`SBC_izy & T==`Tfour & phi2)
			 | (OP==`SBC_izy & T==`Tfive & phi1)
			 | (OP==`SBC_izy & T==`Tfive & phi2)
			 | (OP==`SBC_zpx & T==`Tzero & phi1)
			 | (OP==`SBC_zpx & T==`Tzero & phi2)
			 | (OP==`SBC_zpx & T==`Tone & phi1 & !decMode)
			 | (OP==`SBC_zpx & T==`Tone & phi2 & !decMode)
			 | (OP==`SBC_zpx & T==`Ttwo & phi1)
			 | (OP==`SBC_zpx & T==`Ttwo & phi2)
			 | (OP==`SBC_zpx & T==`Tthree & phi1)
			 | (OP==`SBC_zpx & T==`Tthree & phi2)
			 | (OP==`INC_zpx & T==`Tzero & phi1)
			 | (OP==`INC_zpx & T==`Tzero & phi2)
			 | (OP==`INC_zpx & T==`Tone & phi1)
			 | (OP==`INC_zpx & T==`Tone & phi2)
			 | (OP==`INC_zpx & T==`Ttwo & phi1)
			 | (OP==`INC_zpx & T==`Ttwo & phi2)
			 | (OP==`INC_zpx & T==`Tthree & phi1)
			 | (OP==`INC_zpx & T==`Tthree & phi2)
			 | (OP==`INC_zpx & T==`Tfour & phi1)
			 | (OP==`INC_zpx & T==`Tfour & phi2)
			 | (OP==`INC_zpx & T==`Tfive & phi1)
			 | (OP==`INC_zpx & T==`Tfive & phi2)
			 | (OP==`SED & T==`Tone & phi1)
			 | (OP==`SED & T==`Tone & phi2)
			 | (OP==`SED & T==`Ttwo & phi1)
			 | (OP==`SED & T==`Ttwo & phi2)
			 | (OP==`SBC_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`SBC_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`SBC_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`SBC_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`SBC_aby & T==`Tone & phi1 & !decMode)
			 | (OP==`SBC_aby & T==`Tone & phi2 & !decMode)
			 | (OP==`SBC_aby & T==`Ttwo & phi1)
			 | (OP==`SBC_aby & T==`Ttwo & phi2)
			 | (OP==`SBC_aby & T==`Tthree & phi1)
			 | (OP==`SBC_aby & T==`Tthree & phi2)
			 | (OP==`SBC_aby & T==`Tfour & phi1)
			 | (OP==`SBC_aby & T==`Tfour & phi2)
			 | (OP==`SBC_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`SBC_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`SBC_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`SBC_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`SBC_abx & T==`Tone & phi1 & !decMode)
			 | (OP==`SBC_abx & T==`Tone & phi2 & !decMode)
			 | (OP==`SBC_abx & T==`Ttwo & phi1)
			 | (OP==`SBC_abx & T==`Ttwo & phi2)
			 | (OP==`SBC_abx & T==`Tthree & phi1)
			 | (OP==`SBC_abx & T==`Tthree & phi2)
			 | (OP==`SBC_abx & T==`Tfour & phi1)
			 | (OP==`SBC_abx & T==`Tfour & phi2)
			 | (OP==`INC_abx & T==`Tzero & phi1)
			 | (OP==`INC_abx & T==`Tzero & phi2)
			 | (OP==`INC_abx & T==`Tone & phi1)
			 | (OP==`INC_abx & T==`Tone & phi2)
			 | (OP==`INC_abx & T==`Ttwo & phi1)
			 | (OP==`INC_abx & T==`Ttwo & phi2)
			 | (OP==`INC_abx & T==`Tthree & phi1)
			 | (OP==`INC_abx & T==`Tthree & phi2)
			 | (OP==`INC_abx & T==`Tfour & phi1)
			 | (OP==`INC_abx & T==`Tfour & phi2)
			 | (OP==`INC_abx & T==`Tfive & phi1)
			 | (OP==`INC_abx & T==`Tfive & phi2)
			 | (OP==`INC_abx & T==`Tsix & phi1)
			 | (OP==`INC_abx & T==`Tsix & phi2)
			;

assign control[`SUMS] = (OP==`BRK & T==`Tzero & phi1)
			 | (OP==`BRK & T==`Tzero & phi2)
			 | (OP==`BRK & T==`Tone & phi1)
			 | (OP==`BRK & T==`Tone & phi2)
			 | (OP==`BRK & T==`Ttwo & phi1)
			 | (OP==`BRK & T==`Ttwo & phi2)
			 | (OP==`BRK & T==`Tthree & phi1)
			 | (OP==`BRK & T==`Tthree & phi2)
			 | (OP==`BRK & T==`Tfour & phi1)
			 | (OP==`BRK & T==`Tfour & phi2)
			 | (OP==`BRK & T==`Tfive & phi1)
			 | (OP==`BRK & T==`Tfive & phi2)
			 | (OP==`BRK & T==`Tsix & phi1)
			 | (OP==`BRK & T==`Tsix & phi2)
			 | (OP==`ORA_izx & T==`Tzero & phi1)
			 | (OP==`ORA_izx & T==`Tzero & phi2)
			 | (OP==`ORA_izx & T==`Ttwo & phi1)
			 | (OP==`ORA_izx & T==`Ttwo & phi2)
			 | (OP==`ORA_izx & T==`Tthree & phi1)
			 | (OP==`ORA_izx & T==`Tthree & phi2)
			 | (OP==`ORA_izx & T==`Tfour & phi1)
			 | (OP==`ORA_izx & T==`Tfour & phi2)
			 | (OP==`ORA_izx & T==`Tfive & phi1)
			 | (OP==`ORA_izx & T==`Tfive & phi2)
			 | (OP==`ORA_zp & T==`Tzero & phi1)
			 | (OP==`ORA_zp & T==`Tzero & phi2)
			 | (OP==`ORA_zp & T==`Ttwo & phi1)
			 | (OP==`ORA_zp & T==`Ttwo & phi2)
			 | (OP==`ASL_zp & T==`Tzero & phi1)
			 | (OP==`ASL_zp & T==`Tzero & phi2)
			 | (OP==`ASL_zp & T==`Tone & phi1)
			 | (OP==`ASL_zp & T==`Tone & phi2)
			 | (OP==`ASL_zp & T==`Ttwo & phi1)
			 | (OP==`ASL_zp & T==`Ttwo & phi2)
			 | (OP==`ASL_zp & T==`Tthree & phi1)
			 | (OP==`ASL_zp & T==`Tthree & phi2)
			 | (OP==`ASL_zp & T==`Tfour & phi1)
			 | (OP==`ASL_zp & T==`Tfour & phi2)
			 | (OP==`PHP & T==`Tzero & phi1)
			 | (OP==`PHP & T==`Tzero & phi2)
			 | (OP==`PHP & T==`Tone & phi1)
			 | (OP==`PHP & T==`Tone & phi2)
			 | (OP==`PHP & T==`Ttwo & phi1)
			 | (OP==`PHP & T==`Ttwo & phi2)
			 | (OP==`ORA_imm & T==`Ttwo & phi1)
			 | (OP==`ORA_imm & T==`Ttwo & phi2)
			 | (OP==`ASL & T==`Tone & phi1)
			 | (OP==`ASL & T==`Tone & phi2)
			 | (OP==`ASL & T==`Ttwo & phi1)
			 | (OP==`ASL & T==`Ttwo & phi2)
			 | (OP==`ORA_abs & T==`Tzero & phi1)
			 | (OP==`ORA_abs & T==`Tzero & phi2)
			 | (OP==`ORA_abs & T==`Ttwo & phi1)
			 | (OP==`ORA_abs & T==`Ttwo & phi2)
			 | (OP==`ORA_abs & T==`Tthree & phi1)
			 | (OP==`ORA_abs & T==`Tthree & phi2)
			 | (OP==`ASL_abs & T==`Tzero & phi1)
			 | (OP==`ASL_abs & T==`Tzero & phi2)
			 | (OP==`ASL_abs & T==`Tone & phi1)
			 | (OP==`ASL_abs & T==`Ttwo & phi1)
			 | (OP==`ASL_abs & T==`Ttwo & phi2)
			 | (OP==`ASL_abs & T==`Tthree & phi1)
			 | (OP==`ASL_abs & T==`Tthree & phi2)
			 | (OP==`ASL_abs & T==`Tfour & phi1)
			 | (OP==`ASL_abs & T==`Tfour & phi2)
			 | (OP==`ASL_abs & T==`Tfive & phi1)
			 | (OP==`ASL_abs & T==`Tfive & phi2)
			 | (OP==`BPL_rel & T==`Tzero & phi1)
			 | (OP==`BPL_rel & T==`Tzero & phi2)
			 | (OP==`BPL_rel & T==`Ttwo & phi1)
			 | (OP==`BPL_rel & T==`Ttwo & phi2)
			 | (OP==`BPL_rel & T==`Tthree & phi1)
			 | (OP==`BPL_rel & T==`Tthree & phi2)
			 | (OP==`BPL_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BPL_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BPL_rel & T==`T1BranchCross & phi1)
			 | (OP==`BPL_rel & T==`T1BranchCross & phi2)
			 | (OP==`BPL_rel & T==`T1NoBranch & phi1)
			 | (OP==`BPL_rel & T==`T1NoBranch & phi2)
			 | (OP==`ORA_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`ORA_izy & T==`TzeroCrossPg & phi2)
			 | (OP==`ORA_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ORA_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`ORA_izy & T==`Ttwo & phi1)
			 | (OP==`ORA_izy & T==`Ttwo & phi2)
			 | (OP==`ORA_izy & T==`Tthree & phi1)
			 | (OP==`ORA_izy & T==`Tthree & phi2)
			 | (OP==`ORA_izy & T==`Tfour & phi1)
			 | (OP==`ORA_izy & T==`Tfour & phi2)
			 | (OP==`ORA_izy & T==`Tfive & phi1)
			 | (OP==`ORA_izy & T==`Tfive & phi2)
			 | (OP==`ORA_zpx & T==`Tzero & phi1)
			 | (OP==`ORA_zpx & T==`Tzero & phi2)
			 | (OP==`ORA_zpx & T==`Ttwo & phi1)
			 | (OP==`ORA_zpx & T==`Ttwo & phi2)
			 | (OP==`ORA_zpx & T==`Tthree & phi1)
			 | (OP==`ORA_zpx & T==`Tthree & phi2)
			 | (OP==`ASL_zpx & T==`Tzero & phi1)
			 | (OP==`ASL_zpx & T==`Tzero & phi2)
			 | (OP==`ASL_zpx & T==`Tone & phi1)
			 | (OP==`ASL_zpx & T==`Tone & phi2)
			 | (OP==`ASL_zpx & T==`Ttwo & phi1)
			 | (OP==`ASL_zpx & T==`Ttwo & phi2)
			 | (OP==`ASL_zpx & T==`Tthree & phi1)
			 | (OP==`ASL_zpx & T==`Tthree & phi2)
			 | (OP==`ASL_zpx & T==`Tfour & phi1)
			 | (OP==`ASL_zpx & T==`Tfour & phi2)
			 | (OP==`ASL_zpx & T==`Tfive & phi1)
			 | (OP==`ASL_zpx & T==`Tfive & phi2)
			 | (OP==`CLC & T==`Tone & phi1)
			 | (OP==`CLC & T==`Tone & phi2)
			 | (OP==`CLC & T==`Ttwo & phi1)
			 | (OP==`CLC & T==`Ttwo & phi2)
			 | (OP==`ORA_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ORA_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`ORA_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`ORA_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`ORA_aby & T==`Ttwo & phi1)
			 | (OP==`ORA_aby & T==`Ttwo & phi2)
			 | (OP==`ORA_aby & T==`Tthree & phi1)
			 | (OP==`ORA_aby & T==`Tthree & phi2)
			 | (OP==`ORA_aby & T==`Tfour & phi1)
			 | (OP==`ORA_aby & T==`Tfour & phi2)
			 | (OP==`ORA_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ORA_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`ORA_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`ORA_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`ORA_abx & T==`Ttwo & phi1)
			 | (OP==`ORA_abx & T==`Ttwo & phi2)
			 | (OP==`ORA_abx & T==`Tthree & phi1)
			 | (OP==`ORA_abx & T==`Tthree & phi2)
			 | (OP==`ORA_abx & T==`Tfour & phi1)
			 | (OP==`ORA_abx & T==`Tfour & phi2)
			 | (OP==`ASL_abx & T==`Tzero & phi1)
			 | (OP==`ASL_abx & T==`Tzero & phi2)
			 | (OP==`ASL_abx & T==`Tone & phi1)
			 | (OP==`ASL_abx & T==`Tone & phi2)
			 | (OP==`ASL_abx & T==`Ttwo & phi1)
			 | (OP==`ASL_abx & T==`Ttwo & phi2)
			 | (OP==`ASL_abx & T==`Tthree & phi1)
			 | (OP==`ASL_abx & T==`Tthree & phi2)
			 | (OP==`ASL_abx & T==`Tfour & phi1)
			 | (OP==`ASL_abx & T==`Tfour & phi2)
			 | (OP==`ASL_abx & T==`Tfive & phi1)
			 | (OP==`ASL_abx & T==`Tfive & phi2)
			 | (OP==`ASL_abx & T==`Tsix & phi1)
			 | (OP==`ASL_abx & T==`Tsix & phi2)
			 | (OP==`JSR_abs & T==`Tzero & phi1)
			 | (OP==`JSR_abs & T==`Tzero & phi2)
			 | (OP==`JSR_abs & T==`Tone & phi1)
			 | (OP==`JSR_abs & T==`Tone & phi2)
			 | (OP==`JSR_abs & T==`Ttwo & phi1)
			 | (OP==`JSR_abs & T==`Ttwo & phi2)
			 | (OP==`JSR_abs & T==`Tthree & phi1)
			 | (OP==`JSR_abs & T==`Tthree & phi2)
			 | (OP==`JSR_abs & T==`Tfour & phi1)
			 | (OP==`JSR_abs & T==`Tfour & phi2)
			 | (OP==`JSR_abs & T==`Tfive & phi1)
			 | (OP==`JSR_abs & T==`Tfive & phi2)
			 | (OP==`AND_izx & T==`Tzero & phi1)
			 | (OP==`AND_izx & T==`Tzero & phi2)
			 | (OP==`AND_izx & T==`Ttwo & phi1)
			 | (OP==`AND_izx & T==`Ttwo & phi2)
			 | (OP==`AND_izx & T==`Tthree & phi1)
			 | (OP==`AND_izx & T==`Tthree & phi2)
			 | (OP==`AND_izx & T==`Tfour & phi1)
			 | (OP==`AND_izx & T==`Tfour & phi2)
			 | (OP==`AND_izx & T==`Tfive & phi1)
			 | (OP==`AND_izx & T==`Tfive & phi2)
			 | (OP==`BIT_zp & T==`Tzero & phi1)
			 | (OP==`BIT_zp & T==`Tzero & phi2)
			 | (OP==`BIT_zp & T==`Ttwo & phi1)
			 | (OP==`BIT_zp & T==`Ttwo & phi2)
			 | (OP==`AND_zp & T==`Tzero & phi1)
			 | (OP==`AND_zp & T==`Tzero & phi2)
			 | (OP==`AND_zp & T==`Ttwo & phi1)
			 | (OP==`AND_zp & T==`Ttwo & phi2)
			 | (OP==`ROL_zp & T==`Tzero & phi1)
			 | (OP==`ROL_zp & T==`Tzero & phi2)
			 | (OP==`ROL_zp & T==`Tone & phi1)
			 | (OP==`ROL_zp & T==`Tone & phi2)
			 | (OP==`ROL_zp & T==`Ttwo & phi1)
			 | (OP==`ROL_zp & T==`Ttwo & phi2)
			 | (OP==`ROL_zp & T==`Tthree & phi1)
			 | (OP==`ROL_zp & T==`Tthree & phi2)
			 | (OP==`ROL_zp & T==`Tfour & phi1)
			 | (OP==`ROL_zp & T==`Tfour & phi2)
			 | (OP==`PLP & T==`Tzero & phi1)
			 | (OP==`PLP & T==`Tzero & phi2)
			 | (OP==`PLP & T==`Tone & phi1)
			 | (OP==`PLP & T==`Tone & phi2)
			 | (OP==`PLP & T==`Ttwo & phi1)
			 | (OP==`PLP & T==`Ttwo & phi2)
			 | (OP==`PLP & T==`Tthree & phi1)
			 | (OP==`PLP & T==`Tthree & phi2)
			 | (OP==`AND_imm & T==`Ttwo & phi1)
			 | (OP==`AND_imm & T==`Ttwo & phi2)
			 | (OP==`ROL & T==`Tone & phi1)
			 | (OP==`ROL & T==`Tone & phi2)
			 | (OP==`ROL & T==`Ttwo & phi1)
			 | (OP==`ROL & T==`Ttwo & phi2)
			 | (OP==`BIT_abs & T==`Tzero & phi1)
			 | (OP==`BIT_abs & T==`Tzero & phi2)
			 | (OP==`BIT_abs & T==`Ttwo & phi1)
			 | (OP==`BIT_abs & T==`Ttwo & phi2)
			 | (OP==`BIT_abs & T==`Tthree & phi1)
			 | (OP==`BIT_abs & T==`Tthree & phi2)
			 | (OP==`AND_abs & T==`Tzero & phi1)
			 | (OP==`AND_abs & T==`Tzero & phi2)
			 | (OP==`AND_abs & T==`Ttwo & phi1)
			 | (OP==`AND_abs & T==`Ttwo & phi2)
			 | (OP==`AND_abs & T==`Tthree & phi1)
			 | (OP==`AND_abs & T==`Tthree & phi2)
			 | (OP==`ROL_abs & T==`Tzero & phi1)
			 | (OP==`ROL_abs & T==`Tzero & phi2)
			 | (OP==`ROL_abs & T==`Tone & phi1)
			 | (OP==`ROL_abs & T==`Tone & phi2)
			 | (OP==`ROL_abs & T==`Ttwo & phi1)
			 | (OP==`ROL_abs & T==`Ttwo & phi2)
			 | (OP==`ROL_abs & T==`Tthree & phi1)
			 | (OP==`ROL_abs & T==`Tthree & phi2)
			 | (OP==`ROL_abs & T==`Tfour & phi1)
			 | (OP==`ROL_abs & T==`Tfour & phi2)
			 | (OP==`ROL_abs & T==`Tfive & phi1)
			 | (OP==`ROL_abs & T==`Tfive & phi2)
			 | (OP==`BMI_rel & T==`Tzero & phi1)
			 | (OP==`BMI_rel & T==`Tzero & phi2)
			 | (OP==`BMI_rel & T==`Ttwo & phi1)
			 | (OP==`BMI_rel & T==`Ttwo & phi2)
			 | (OP==`BMI_rel & T==`Tthree & phi1)
			 | (OP==`BMI_rel & T==`Tthree & phi2)
			 | (OP==`BMI_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BMI_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BMI_rel & T==`T1BranchCross & phi1)
			 | (OP==`BMI_rel & T==`T1BranchCross & phi2)
			 | (OP==`BMI_rel & T==`T1NoBranch & phi1)
			 | (OP==`BMI_rel & T==`T1NoBranch & phi2)
			 | (OP==`AND_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`AND_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`AND_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`AND_izy & T==`TzeroCrossPg & phi2)
			 | (OP==`AND_izy & T==`Ttwo & phi1)
			 | (OP==`AND_izy & T==`Ttwo & phi2)
			 | (OP==`AND_izy & T==`Tthree & phi1)
			 | (OP==`AND_izy & T==`Tthree & phi2)
			 | (OP==`AND_izy & T==`Tfour & phi1)
			 | (OP==`AND_izy & T==`Tfour & phi2)
			 | (OP==`AND_izy & T==`Tfive & phi1)
			 | (OP==`AND_izy & T==`Tfive & phi2)
			 | (OP==`AND_zpx & T==`Tzero & phi1)
			 | (OP==`AND_zpx & T==`Tzero & phi2)
			 | (OP==`AND_zpx & T==`Ttwo & phi1)
			 | (OP==`AND_zpx & T==`Ttwo & phi2)
			 | (OP==`AND_zpx & T==`Tthree & phi1)
			 | (OP==`AND_zpx & T==`Tthree & phi2)
			 | (OP==`ROL_zpx & T==`Tzero & phi1)
			 | (OP==`ROL_zpx & T==`Tzero & phi2)
			 | (OP==`ROL_zpx & T==`Tone & phi1)
			 | (OP==`ROL_zpx & T==`Tone & phi2)
			 | (OP==`ROL_zpx & T==`Ttwo & phi1)
			 | (OP==`ROL_zpx & T==`Ttwo & phi2)
			 | (OP==`ROL_zpx & T==`Tthree & phi1)
			 | (OP==`ROL_zpx & T==`Tthree & phi2)
			 | (OP==`ROL_zpx & T==`Tfour & phi1)
			 | (OP==`ROL_zpx & T==`Tfour & phi2)
			 | (OP==`ROL_zpx & T==`Tfive & phi1)
			 | (OP==`ROL_zpx & T==`Tfive & phi2)
			 | (OP==`SEC & T==`Tone & phi1)
			 | (OP==`SEC & T==`Tone & phi2)
			 | (OP==`SEC & T==`Ttwo & phi1)
			 | (OP==`SEC & T==`Ttwo & phi2)
			 | (OP==`AND_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`AND_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`AND_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`AND_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`AND_aby & T==`Ttwo & phi1)
			 | (OP==`AND_aby & T==`Ttwo & phi2)
			 | (OP==`AND_aby & T==`Tthree & phi1)
			 | (OP==`AND_aby & T==`Tthree & phi2)
			 | (OP==`AND_aby & T==`Tfour & phi1)
			 | (OP==`AND_aby & T==`Tfour & phi2)
			 | (OP==`AND_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`AND_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`AND_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`AND_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`AND_abx & T==`Ttwo & phi1)
			 | (OP==`AND_abx & T==`Ttwo & phi2)
			 | (OP==`AND_abx & T==`Tthree & phi1)
			 | (OP==`AND_abx & T==`Tthree & phi2)
			 | (OP==`AND_abx & T==`Tfour & phi1)
			 | (OP==`AND_abx & T==`Tfour & phi2)
			 | (OP==`ROL_abx & T==`Tzero & phi1)
			 | (OP==`ROL_abx & T==`Tzero & phi2)
			 | (OP==`ROL_abx & T==`Tone & phi1)
			 | (OP==`ROL_abx & T==`Tone & phi2)
			 | (OP==`ROL_abx & T==`Ttwo & phi1)
			 | (OP==`ROL_abx & T==`Ttwo & phi2)
			 | (OP==`ROL_abx & T==`Tthree & phi1)
			 | (OP==`ROL_abx & T==`Tthree & phi2)
			 | (OP==`ROL_abx & T==`Tfour & phi1)
			 | (OP==`ROL_abx & T==`Tfour & phi2)
			 | (OP==`ROL_abx & T==`Tfive & phi1)
			 | (OP==`ROL_abx & T==`Tfive & phi2)
			 | (OP==`ROL_abx & T==`Tsix & phi1)
			 | (OP==`ROL_abx & T==`Tsix & phi2)
			 | (OP==`RTI & T==`Tzero & phi1)
			 | (OP==`RTI & T==`Tzero & phi2)
			 | (OP==`RTI & T==`Tone & phi1)
			 | (OP==`RTI & T==`Tone & phi2)
			 | (OP==`RTI & T==`Ttwo & phi1)
			 | (OP==`RTI & T==`Ttwo & phi2)
			 | (OP==`RTI & T==`Tthree & phi1)
			 | (OP==`RTI & T==`Tthree & phi2)
			 | (OP==`RTI & T==`Tfour & phi1)
			 | (OP==`RTI & T==`Tfour & phi2)
			 | (OP==`RTI & T==`Tfive & phi1)
			 | (OP==`RTI & T==`Tfive & phi2)
			 | (OP==`EOR_izx & T==`Tzero & phi1)
			 | (OP==`EOR_izx & T==`Tzero & phi2)
			 | (OP==`EOR_izx & T==`Ttwo & phi1)
			 | (OP==`EOR_izx & T==`Ttwo & phi2)
			 | (OP==`EOR_izx & T==`Tthree & phi1)
			 | (OP==`EOR_izx & T==`Tthree & phi2)
			 | (OP==`EOR_izx & T==`Tfour & phi1)
			 | (OP==`EOR_izx & T==`Tfour & phi2)
			 | (OP==`EOR_izx & T==`Tfive & phi1)
			 | (OP==`EOR_izx & T==`Tfive & phi2)
			 | (OP==`EOR_zp & T==`Tzero & phi1)
			 | (OP==`EOR_zp & T==`Tzero & phi2)
			 | (OP==`EOR_zp & T==`Ttwo & phi1)
			 | (OP==`EOR_zp & T==`Ttwo & phi2)
			 | (OP==`LSR_zp & T==`Tzero & phi1)
			 | (OP==`LSR_zp & T==`Tzero & phi2)
			 | (OP==`LSR_zp & T==`Tone & phi1)
			 | (OP==`LSR_zp & T==`Tone & phi2)
			 | (OP==`LSR_zp & T==`Ttwo & phi1)
			 | (OP==`LSR_zp & T==`Ttwo & phi2)
			 | (OP==`LSR_zp & T==`Tthree & phi1)
			 | (OP==`LSR_zp & T==`Tthree & phi2)
			 | (OP==`PHA & T==`Tzero & phi1)
			 | (OP==`PHA & T==`Tzero & phi2)
			 | (OP==`PHA & T==`Tone & phi1)
			 | (OP==`PHA & T==`Tone & phi2)
			 | (OP==`PHA & T==`Ttwo & phi1)
			 | (OP==`PHA & T==`Ttwo & phi2)
			 | (OP==`EOR_imm & T==`Ttwo & phi1)
			 | (OP==`EOR_imm & T==`Ttwo & phi2)
			 | (OP==`LSR & T==`Ttwo & phi1)
			 | (OP==`LSR & T==`Ttwo & phi2)
			 | (OP==`JMP_abs & T==`Tzero & phi1)
			 | (OP==`JMP_abs & T==`Tzero & phi2)
			 | (OP==`JMP_abs & T==`Tone & phi1)
			 | (OP==`JMP_abs & T==`Tone & phi2)
			 | (OP==`JMP_abs & T==`Ttwo & phi1)
			 | (OP==`JMP_abs & T==`Ttwo & phi2)
			 | (OP==`EOR_abs & T==`Tzero & phi1)
			 | (OP==`EOR_abs & T==`Tzero & phi2)
			 | (OP==`EOR_abs & T==`Ttwo & phi1)
			 | (OP==`EOR_abs & T==`Ttwo & phi2)
			 | (OP==`EOR_abs & T==`Tthree & phi1)
			 | (OP==`EOR_abs & T==`Tthree & phi2)
			 | (OP==`LSR_abs & T==`Tzero & phi1)
			 | (OP==`LSR_abs & T==`Tzero & phi2)
			 | (OP==`LSR_abs & T==`Tone & phi1)
			 | (OP==`LSR_abs & T==`Tone & phi2)
			 | (OP==`LSR_abs & T==`Ttwo & phi1)
			 | (OP==`LSR_abs & T==`Ttwo & phi2)
			 | (OP==`LSR_abs & T==`Tthree & phi1)
			 | (OP==`LSR_abs & T==`Tthree & phi2)
			 | (OP==`LSR_abs & T==`Tfour & phi1)
			 | (OP==`LSR_abs & T==`Tfour & phi2)
			 | (OP==`BVC_rel & T==`Tzero & phi1)
			 | (OP==`BVC_rel & T==`Tzero & phi2)
			 | (OP==`BVC_rel & T==`Ttwo & phi1)
			 | (OP==`BVC_rel & T==`Ttwo & phi2)
			 | (OP==`BVC_rel & T==`Tthree & phi1)
			 | (OP==`BVC_rel & T==`Tthree & phi2)
			 | (OP==`BVC_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BVC_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BVC_rel & T==`T1BranchCross & phi1)
			 | (OP==`BVC_rel & T==`T1BranchCross & phi2)
			 | (OP==`BVC_rel & T==`T1NoBranch & phi1)
			 | (OP==`BVC_rel & T==`T1NoBranch & phi2)
			 | (OP==`EOR_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`EOR_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`EOR_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`EOR_izy & T==`TzeroCrossPg & phi2)
			 | (OP==`EOR_izy & T==`Ttwo & phi1)
			 | (OP==`EOR_izy & T==`Ttwo & phi2)
			 | (OP==`EOR_izy & T==`Tthree & phi1)
			 | (OP==`EOR_izy & T==`Tthree & phi2)
			 | (OP==`EOR_izy & T==`Tfour & phi1)
			 | (OP==`EOR_izy & T==`Tfour & phi2)
			 | (OP==`EOR_izy & T==`Tfive & phi1)
			 | (OP==`EOR_izy & T==`Tfive & phi2)
			 | (OP==`EOR_zpx & T==`Tzero & phi1)
			 | (OP==`EOR_zpx & T==`Tzero & phi2)
			 | (OP==`EOR_zpx & T==`Ttwo & phi1)
			 | (OP==`EOR_zpx & T==`Ttwo & phi2)
			 | (OP==`EOR_zpx & T==`Tthree & phi1)
			 | (OP==`EOR_zpx & T==`Tthree & phi2)
			 | (OP==`LSR_zpx & T==`Tzero & phi1)
			 | (OP==`LSR_zpx & T==`Tzero & phi2)
			 | (OP==`LSR_zpx & T==`Tone & phi1)
			 | (OP==`LSR_zpx & T==`Tone & phi2)
			 | (OP==`LSR_zpx & T==`Ttwo & phi1)
			 | (OP==`LSR_zpx & T==`Ttwo & phi2)
			 | (OP==`LSR_zpx & T==`Tthree & phi1)
			 | (OP==`LSR_zpx & T==`Tthree & phi2)
			 | (OP==`LSR_zpx & T==`Tfour & phi1)
			 | (OP==`LSR_zpx & T==`Tfour & phi2)
			 | (OP==`CLI & T==`Tone & phi1)
			 | (OP==`CLI & T==`Tone & phi2)
			 | (OP==`CLI & T==`Ttwo & phi1)
			 | (OP==`CLI & T==`Ttwo & phi2)
			 | (OP==`EOR_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`EOR_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`EOR_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`EOR_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`EOR_aby & T==`Ttwo & phi1)
			 | (OP==`EOR_aby & T==`Ttwo & phi2)
			 | (OP==`EOR_aby & T==`Tthree & phi1)
			 | (OP==`EOR_aby & T==`Tthree & phi2)
			 | (OP==`EOR_aby & T==`Tfour & phi1)
			 | (OP==`EOR_aby & T==`Tfour & phi2)
			 | (OP==`EOR_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`EOR_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`EOR_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`EOR_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`EOR_abx & T==`Ttwo & phi1)
			 | (OP==`EOR_abx & T==`Ttwo & phi2)
			 | (OP==`EOR_abx & T==`Tthree & phi1)
			 | (OP==`EOR_abx & T==`Tthree & phi2)
			 | (OP==`EOR_abx & T==`Tfour & phi1)
			 | (OP==`EOR_abx & T==`Tfour & phi2)
			 | (OP==`LSR_abx & T==`Tzero & phi1)
			 | (OP==`LSR_abx & T==`Tzero & phi2)
			 | (OP==`LSR_abx & T==`Tone & phi1)
			 | (OP==`LSR_abx & T==`Tone & phi2)
			 | (OP==`LSR_abx & T==`Ttwo & phi1)
			 | (OP==`LSR_abx & T==`Ttwo & phi2)
			 | (OP==`LSR_abx & T==`Tthree & phi1)
			 | (OP==`LSR_abx & T==`Tthree & phi2)
			 | (OP==`LSR_abx & T==`Tfour & phi1)
			 | (OP==`LSR_abx & T==`Tfour & phi2)
			 | (OP==`LSR_abx & T==`Tfive & phi1)
			 | (OP==`LSR_abx & T==`Tfive & phi2)
			 | (OP==`RTS & T==`Tzero & phi1)
			 | (OP==`RTS & T==`Tzero & phi2)
			 | (OP==`RTS & T==`Tone & phi1)
			 | (OP==`RTS & T==`Tone & phi2)
			 | (OP==`RTS & T==`Ttwo & phi1)
			 | (OP==`RTS & T==`Ttwo & phi2)
			 | (OP==`RTS & T==`Tthree & phi1)
			 | (OP==`RTS & T==`Tthree & phi2)
			 | (OP==`RTS & T==`Tfour & phi1)
			 | (OP==`RTS & T==`Tfour & phi2)
			 | (OP==`RTS & T==`Tfive & phi1)
			 | (OP==`RTS & T==`Tfive & phi2)
			 | (OP==`ADC_izx & T==`Tzero & phi1)
			 | (OP==`ADC_izx & T==`Tzero & phi2)
			 | (OP==`ADC_izx & T==`Tone & phi1)
			 | (OP==`ADC_izx & T==`Tone & phi2)
			 | (OP==`ADC_izx & T==`Ttwo & phi1)
			 | (OP==`ADC_izx & T==`Ttwo & phi2)
			 | (OP==`ADC_izx & T==`Tthree & phi1)
			 | (OP==`ADC_izx & T==`Tthree & phi2)
			 | (OP==`ADC_izx & T==`Tfour & phi1)
			 | (OP==`ADC_izx & T==`Tfour & phi2)
			 | (OP==`ADC_izx & T==`Tfive & phi1)
			 | (OP==`ADC_izx & T==`Tfive & phi2)
			 | (OP==`ADC_zp & T==`Tzero & phi1)
			 | (OP==`ADC_zp & T==`Tzero & phi2)
			 | (OP==`ADC_zp & T==`Tone & phi1)
			 | (OP==`ADC_zp & T==`Tone & phi2)
			 | (OP==`ADC_zp & T==`Ttwo & phi1)
			 | (OP==`ADC_zp & T==`Ttwo & phi2)
			 | (OP==`ROR_zp & T==`Tzero & phi1)
			 | (OP==`ROR_zp & T==`Tzero & phi2)
			 | (OP==`ROR_zp & T==`Tone & phi1)
			 | (OP==`ROR_zp & T==`Tone & phi2)
			 | (OP==`ROR_zp & T==`Ttwo & phi1)
			 | (OP==`ROR_zp & T==`Ttwo & phi2)
			 | (OP==`ROR_zp & T==`Tthree & phi1)
			 | (OP==`ROR_zp & T==`Tthree & phi2)
			 | (OP==`PLA & T==`Tzero & phi1)
			 | (OP==`PLA & T==`Tzero & phi2)
			 | (OP==`PLA & T==`Tone & phi1)
			 | (OP==`PLA & T==`Tone & phi2)
			 | (OP==`PLA & T==`Ttwo & phi1)
			 | (OP==`PLA & T==`Ttwo & phi2)
			 | (OP==`PLA & T==`Tthree & phi1)
			 | (OP==`PLA & T==`Tthree & phi2)
			 | (OP==`ADC_imm & T==`Tone & phi1)
			 | (OP==`ADC_imm & T==`Tone & phi2)
			 | (OP==`ADC_imm & T==`Ttwo & phi1)
			 | (OP==`ADC_imm & T==`Ttwo & phi2)
			 | (OP==`ROR & T==`Ttwo & phi1)
			 | (OP==`ROR & T==`Ttwo & phi2)
			 | (OP==`JMP_zp & T==`Tzero & phi1)
			 | (OP==`JMP_zp & T==`Tzero & phi2)
			 | (OP==`JMP_zp & T==`Tone & phi1)
			 | (OP==`JMP_zp & T==`Tone & phi2)
			 | (OP==`JMP_zp & T==`Ttwo & phi1)
			 | (OP==`JMP_zp & T==`Ttwo & phi2)
			 | (OP==`JMP_zp & T==`Tthree & phi1)
			 | (OP==`JMP_zp & T==`Tthree & phi2)
			 | (OP==`JMP_zp & T==`Tfour & phi1)
			 | (OP==`JMP_zp & T==`Tfour & phi2)
			 | (OP==`ADC_abs & T==`Tzero & phi1)
			 | (OP==`ADC_abs & T==`Tzero & phi2)
			 | (OP==`ADC_abs & T==`Tone & phi1)
			 | (OP==`ADC_abs & T==`Tone & phi2)
			 | (OP==`ADC_abs & T==`Ttwo & phi1)
			 | (OP==`ADC_abs & T==`Ttwo & phi2)
			 | (OP==`ADC_abs & T==`Tthree & phi1)
			 | (OP==`ADC_abs & T==`Tthree & phi2)
			 | (OP==`ROR_abs & T==`Tzero & phi1)
			 | (OP==`ROR_abs & T==`Tzero & phi2)
			 | (OP==`ROR_abs & T==`Tone & phi1)
			 | (OP==`ROR_abs & T==`Tone & phi2)
			 | (OP==`ROR_abs & T==`Ttwo & phi1)
			 | (OP==`ROR_abs & T==`Ttwo & phi2)
			 | (OP==`ROR_abs & T==`Tthree & phi1)
			 | (OP==`ROR_abs & T==`Tthree & phi2)
			 | (OP==`ROR_abs & T==`Tfour & phi1)
			 | (OP==`ROR_abs & T==`Tfour & phi2)
			 | (OP==`BVS_rel & T==`Tzero & phi1)
			 | (OP==`BVS_rel & T==`Tzero & phi2)
			 | (OP==`BVS_rel & T==`Ttwo & phi1)
			 | (OP==`BVS_rel & T==`Ttwo & phi2)
			 | (OP==`BVS_rel & T==`Tthree & phi1)
			 | (OP==`BVS_rel & T==`Tthree & phi2)
			 | (OP==`BVS_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BVS_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BVS_rel & T==`T1BranchCross & phi1)
			 | (OP==`BVS_rel & T==`T1BranchCross & phi2)
			 | (OP==`BVS_rel & T==`T1NoBranch & phi1)
			 | (OP==`BVS_rel & T==`T1NoBranch & phi2)
			 | (OP==`ADC_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ADC_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`ADC_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`ADC_izy & T==`TzeroCrossPg & phi2)
			 | (OP==`ADC_izy & T==`Tone & phi1)
			 | (OP==`ADC_izy & T==`Tone & phi2)
			 | (OP==`ADC_izy & T==`Ttwo & phi1)
			 | (OP==`ADC_izy & T==`Ttwo & phi2)
			 | (OP==`ADC_izy & T==`Tthree & phi1)
			 | (OP==`ADC_izy & T==`Tthree & phi2)
			 | (OP==`ADC_izy & T==`Tfour & phi1)
			 | (OP==`ADC_izy & T==`Tfour & phi2)
			 | (OP==`ADC_izy & T==`Tfive & phi1)
			 | (OP==`ADC_izy & T==`Tfive & phi2)
			 | (OP==`ADC_zpx & T==`Tzero & phi1)
			 | (OP==`ADC_zpx & T==`Tzero & phi2)
			 | (OP==`ADC_zpx & T==`Tone & phi1)
			 | (OP==`ADC_zpx & T==`Tone & phi2)
			 | (OP==`ADC_zpx & T==`Ttwo & phi1)
			 | (OP==`ADC_zpx & T==`Ttwo & phi2)
			 | (OP==`ADC_zpx & T==`Tthree & phi1)
			 | (OP==`ADC_zpx & T==`Tthree & phi2)
			 | (OP==`ROR_zpx & T==`Tzero & phi1)
			 | (OP==`ROR_zpx & T==`Tzero & phi2)
			 | (OP==`ROR_zpx & T==`Tone & phi1)
			 | (OP==`ROR_zpx & T==`Tone & phi2)
			 | (OP==`ROR_zpx & T==`Ttwo & phi1)
			 | (OP==`ROR_zpx & T==`Ttwo & phi2)
			 | (OP==`ROR_zpx & T==`Tthree & phi1)
			 | (OP==`ROR_zpx & T==`Tthree & phi2)
			 | (OP==`ROR_zpx & T==`Tfour & phi1)
			 | (OP==`ROR_zpx & T==`Tfour & phi2)
			 | (OP==`SEI & T==`Tone & phi1)
			 | (OP==`SEI & T==`Tone & phi2)
			 | (OP==`SEI & T==`Ttwo & phi1)
			 | (OP==`SEI & T==`Ttwo & phi2)
			 | (OP==`ADC_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ADC_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`ADC_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`ADC_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`ADC_aby & T==`Tone & phi1)
			 | (OP==`ADC_aby & T==`Tone & phi2)
			 | (OP==`ADC_aby & T==`Ttwo & phi1)
			 | (OP==`ADC_aby & T==`Ttwo & phi2)
			 | (OP==`ADC_aby & T==`Tthree & phi1)
			 | (OP==`ADC_aby & T==`Tthree & phi2)
			 | (OP==`ADC_aby & T==`Tfour & phi1)
			 | (OP==`ADC_aby & T==`Tfour & phi2)
			 | (OP==`ADC_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ADC_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`ADC_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`ADC_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`ADC_abx & T==`Tone & phi1)
			 | (OP==`ADC_abx & T==`Tone & phi2)
			 | (OP==`ADC_abx & T==`Ttwo & phi1)
			 | (OP==`ADC_abx & T==`Ttwo & phi2)
			 | (OP==`ADC_abx & T==`Tthree & phi1)
			 | (OP==`ADC_abx & T==`Tthree & phi2)
			 | (OP==`ADC_abx & T==`Tfour & phi1)
			 | (OP==`ADC_abx & T==`Tfour & phi2)
			 | (OP==`ROR_abx & T==`Tzero & phi1)
			 | (OP==`ROR_abx & T==`Tzero & phi2)
			 | (OP==`ROR_abx & T==`Tone & phi1)
			 | (OP==`ROR_abx & T==`Tone & phi2)
			 | (OP==`ROR_abx & T==`Ttwo & phi1)
			 | (OP==`ROR_abx & T==`Ttwo & phi2)
			 | (OP==`ROR_abx & T==`Tthree & phi1)
			 | (OP==`ROR_abx & T==`Tthree & phi2)
			 | (OP==`ROR_abx & T==`Tfour & phi1)
			 | (OP==`ROR_abx & T==`Tfour & phi2)
			 | (OP==`ROR_abx & T==`Tfive & phi1)
			 | (OP==`ROR_abx & T==`Tfive & phi2)
			 | (OP==`STA_izx & T==`Tzero & phi1)
			 | (OP==`STA_izx & T==`Tzero & phi2)
			 | (OP==`STA_izx & T==`Tone & phi1)
			 | (OP==`STA_izx & T==`Tone & phi2)
			 | (OP==`STA_izx & T==`Ttwo & phi1)
			 | (OP==`STA_izx & T==`Ttwo & phi2)
			 | (OP==`STA_izx & T==`Tthree & phi1)
			 | (OP==`STA_izx & T==`Tthree & phi2)
			 | (OP==`STA_izx & T==`Tfour & phi1)
			 | (OP==`STA_izx & T==`Tfour & phi2)
			 | (OP==`STA_izx & T==`Tfive & phi1)
			 | (OP==`STA_izx & T==`Tfive & phi2)
			 | (OP==`STY_zp & T==`Tzero & phi1)
			 | (OP==`STY_zp & T==`Tzero & phi2)
			 | (OP==`STY_zp & T==`Tone & phi1)
			 | (OP==`STY_zp & T==`Tone & phi2)
			 | (OP==`STY_zp & T==`Ttwo & phi1)
			 | (OP==`STY_zp & T==`Ttwo & phi2)
			 | (OP==`STA_zp & T==`Tzero & phi1)
			 | (OP==`STA_zp & T==`Tzero & phi2)
			 | (OP==`STA_zp & T==`Tone & phi1)
			 | (OP==`STA_zp & T==`Tone & phi2)
			 | (OP==`STA_zp & T==`Ttwo & phi1)
			 | (OP==`STA_zp & T==`Ttwo & phi2)
			 | (OP==`STX_zp & T==`Tzero & phi1)
			 | (OP==`STX_zp & T==`Tzero & phi2)
			 | (OP==`STX_zp & T==`Tone & phi1)
			 | (OP==`STX_zp & T==`Tone & phi2)
			 | (OP==`STX_zp & T==`Ttwo & phi1)
			 | (OP==`STX_zp & T==`Ttwo & phi2)
			 | (OP==`DEY & T==`Tone & phi1)
			 | (OP==`DEY & T==`Tone & phi2)
			 | (OP==`DEY & T==`Ttwo & phi1)
			 | (OP==`DEY & T==`Ttwo & phi2)
			 | (OP==`TXA & T==`Tone & phi1)
			 | (OP==`TXA & T==`Tone & phi2)
			 | (OP==`TXA & T==`Ttwo & phi1)
			 | (OP==`TXA & T==`Ttwo & phi2)
			 | (OP==`STY_abs & T==`Tzero & phi1)
			 | (OP==`STY_abs & T==`Tzero & phi2)
			 | (OP==`STY_abs & T==`Tone & phi1)
			 | (OP==`STY_abs & T==`Tone & phi2)
			 | (OP==`STY_abs & T==`Ttwo & phi1)
			 | (OP==`STY_abs & T==`Ttwo & phi2)
			 | (OP==`STY_abs & T==`Tthree & phi1)
			 | (OP==`STY_abs & T==`Tthree & phi2)
			 | (OP==`STA_abs & T==`Tzero & phi1)
			 | (OP==`STA_abs & T==`Tzero & phi2)
			 | (OP==`STA_abs & T==`Tone & phi1)
			 | (OP==`STA_abs & T==`Tone & phi2)
			 | (OP==`STA_abs & T==`Ttwo & phi1)
			 | (OP==`STA_abs & T==`Ttwo & phi2)
			 | (OP==`STA_abs & T==`Tthree & phi1)
			 | (OP==`STA_abs & T==`Tthree & phi2)
			 | (OP==`STX_abs & T==`Tzero & phi1)
			 | (OP==`STX_abs & T==`Tzero & phi2)
			 | (OP==`STX_abs & T==`Tone & phi1)
			 | (OP==`STX_abs & T==`Tone & phi2)
			 | (OP==`STX_abs & T==`Ttwo & phi1)
			 | (OP==`STX_abs & T==`Ttwo & phi2)
			 | (OP==`STX_abs & T==`Tthree & phi1)
			 | (OP==`STX_abs & T==`Tthree & phi2)
			 | (OP==`BCC_rel & T==`Tzero & phi1)
			 | (OP==`BCC_rel & T==`Tzero & phi2)
			 | (OP==`BCC_rel & T==`Ttwo & phi1)
			 | (OP==`BCC_rel & T==`Ttwo & phi2)
			 | (OP==`BCC_rel & T==`Tthree & phi1)
			 | (OP==`BCC_rel & T==`Tthree & phi2)
			 | (OP==`BCC_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BCC_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BCC_rel & T==`T1BranchCross & phi1)
			 | (OP==`BCC_rel & T==`T1BranchCross & phi2)
			 | (OP==`BCC_rel & T==`T1NoBranch & phi1)
			 | (OP==`BCC_rel & T==`T1NoBranch & phi2)
			 | (OP==`STA_izy & T==`Tzero & phi1)
			 | (OP==`STA_izy & T==`Tzero & phi2)
			 | (OP==`STA_izy & T==`Tone & phi1)
			 | (OP==`STA_izy & T==`Tone & phi2)
			 | (OP==`STA_izy & T==`Ttwo & phi1)
			 | (OP==`STA_izy & T==`Ttwo & phi2)
			 | (OP==`STA_izy & T==`Tthree & phi1)
			 | (OP==`STA_izy & T==`Tthree & phi2)
			 | (OP==`STA_izy & T==`Tfour & phi1)
			 | (OP==`STA_izy & T==`Tfour & phi2)
			 | (OP==`STA_izy & T==`Tfive & phi1)
			 | (OP==`STA_izy & T==`Tfive & phi2)
			 | (OP==`STY_zpx & T==`Tzero & phi1)
			 | (OP==`STY_zpx & T==`Tzero & phi2)
			 | (OP==`STY_zpx & T==`Tone & phi1)
			 | (OP==`STY_zpx & T==`Tone & phi2)
			 | (OP==`STY_zpx & T==`Ttwo & phi1)
			 | (OP==`STY_zpx & T==`Ttwo & phi2)
			 | (OP==`STY_zpx & T==`Tthree & phi1)
			 | (OP==`STY_zpx & T==`Tthree & phi2)
			 | (OP==`STA_zpx & T==`Tzero & phi1)
			 | (OP==`STA_zpx & T==`Tzero & phi2)
			 | (OP==`STA_zpx & T==`Tone & phi1)
			 | (OP==`STA_zpx & T==`Tone & phi2)
			 | (OP==`STA_zpx & T==`Ttwo & phi1)
			 | (OP==`STA_zpx & T==`Ttwo & phi2)
			 | (OP==`STA_zpx & T==`Tthree & phi1)
			 | (OP==`STA_zpx & T==`Tthree & phi2)
			 | (OP==`STX_zpy & T==`Tzero & phi1)
			 | (OP==`STX_zpy & T==`Tzero & phi2)
			 | (OP==`STX_zpy & T==`Tone & phi1)
			 | (OP==`STX_zpy & T==`Tone & phi2)
			 | (OP==`STX_zpy & T==`Ttwo & phi1)
			 | (OP==`STX_zpy & T==`Ttwo & phi2)
			 | (OP==`STX_zpy & T==`Tthree & phi1)
			 | (OP==`STX_zpy & T==`Tthree & phi2)
			 | (OP==`TYA & T==`Tone & phi1)
			 | (OP==`TYA & T==`Tone & phi2)
			 | (OP==`TYA & T==`Ttwo & phi1)
			 | (OP==`TYA & T==`Ttwo & phi2)
			 | (OP==`STA_aby & T==`Tzero & phi1)
			 | (OP==`STA_aby & T==`Tzero & phi2)
			 | (OP==`STA_aby & T==`Tone & phi1)
			 | (OP==`STA_aby & T==`Tone & phi2)
			 | (OP==`STA_aby & T==`Ttwo & phi1)
			 | (OP==`STA_aby & T==`Ttwo & phi2)
			 | (OP==`STA_aby & T==`Tthree & phi1)
			 | (OP==`STA_aby & T==`Tthree & phi2)
			 | (OP==`STA_aby & T==`Tfour & phi1)
			 | (OP==`STA_aby & T==`Tfour & phi2)
			 | (OP==`TXS & T==`Tone & phi1)
			 | (OP==`TXS & T==`Tone & phi2)
			 | (OP==`TXS & T==`Ttwo & phi1)
			 | (OP==`TXS & T==`Ttwo & phi2)
			 | (OP==`STA_abx & T==`Tzero & phi1)
			 | (OP==`STA_abx & T==`Tzero & phi2)
			 | (OP==`STA_abx & T==`Tone & phi1)
			 | (OP==`STA_abx & T==`Tone & phi2)
			 | (OP==`STA_abx & T==`Ttwo & phi1)
			 | (OP==`STA_abx & T==`Ttwo & phi2)
			 | (OP==`STA_abx & T==`Tthree & phi1)
			 | (OP==`STA_abx & T==`Tthree & phi2)
			 | (OP==`STA_abx & T==`Tfour & phi1)
			 | (OP==`STA_abx & T==`Tfour & phi2)
			 | (OP==`LDY_imm & T==`Tone & phi1)
			 | (OP==`LDY_imm & T==`Tone & phi2)
			 | (OP==`LDY_imm & T==`Ttwo & phi1)
			 | (OP==`LDY_imm & T==`Ttwo & phi2)
			 | (OP==`LDA_izx & T==`Tzero & phi1)
			 | (OP==`LDA_izx & T==`Tzero & phi2)
			 | (OP==`LDA_izx & T==`Tone & phi1)
			 | (OP==`LDA_izx & T==`Tone & phi2)
			 | (OP==`LDA_izx & T==`Ttwo & phi1)
			 | (OP==`LDA_izx & T==`Ttwo & phi2)
			 | (OP==`LDA_izx & T==`Tthree & phi1)
			 | (OP==`LDA_izx & T==`Tthree & phi2)
			 | (OP==`LDA_izx & T==`Tfour & phi1)
			 | (OP==`LDA_izx & T==`Tfour & phi2)
			 | (OP==`LDA_izx & T==`Tfive & phi1)
			 | (OP==`LDA_izx & T==`Tfive & phi2)
			 | (OP==`LDX_imm & T==`Tone & phi1)
			 | (OP==`LDX_imm & T==`Tone & phi2)
			 | (OP==`LDX_imm & T==`Ttwo & phi1)
			 | (OP==`LDX_imm & T==`Ttwo & phi2)
			 | (OP==`LDY_zp & T==`Tzero & phi1)
			 | (OP==`LDY_zp & T==`Tzero & phi2)
			 | (OP==`LDY_zp & T==`Tone & phi1)
			 | (OP==`LDY_zp & T==`Tone & phi2)
			 | (OP==`LDY_zp & T==`Ttwo & phi1)
			 | (OP==`LDY_zp & T==`Ttwo & phi2)
			 | (OP==`LDA_zp & T==`Tzero & phi1)
			 | (OP==`LDA_zp & T==`Tzero & phi2)
			 | (OP==`LDA_zp & T==`Tone & phi1)
			 | (OP==`LDA_zp & T==`Tone & phi2)
			 | (OP==`LDA_zp & T==`Ttwo & phi1)
			 | (OP==`LDA_zp & T==`Ttwo & phi2)
			 | (OP==`LDX_zp & T==`Tzero & phi1)
			 | (OP==`LDX_zp & T==`Tzero & phi2)
			 | (OP==`LDX_zp & T==`Tone & phi1)
			 | (OP==`LDX_zp & T==`Tone & phi2)
			 | (OP==`LDX_zp & T==`Ttwo & phi1)
			 | (OP==`LDX_zp & T==`Ttwo & phi2)
			 | (OP==`TAY & T==`Tone & phi1)
			 | (OP==`TAY & T==`Tone & phi2)
			 | (OP==`TAY & T==`Ttwo & phi1)
			 | (OP==`TAY & T==`Ttwo & phi2)
			 | (OP==`LDA_imm & T==`Tone & phi1)
			 | (OP==`LDA_imm & T==`Tone & phi2)
			 | (OP==`LDA_imm & T==`Ttwo & phi1)
			 | (OP==`LDA_imm & T==`Ttwo & phi2)
			 | (OP==`TAX & T==`Tone & phi1)
			 | (OP==`TAX & T==`Tone & phi2)
			 | (OP==`TAX & T==`Ttwo & phi1)
			 | (OP==`TAX & T==`Ttwo & phi2)
			 | (OP==`LDY_abs & T==`Tzero & phi1)
			 | (OP==`LDY_abs & T==`Tzero & phi2)
			 | (OP==`LDY_abs & T==`Tone & phi1)
			 | (OP==`LDY_abs & T==`Tone & phi2)
			 | (OP==`LDY_abs & T==`Ttwo & phi1)
			 | (OP==`LDY_abs & T==`Ttwo & phi2)
			 | (OP==`LDY_abs & T==`Tthree & phi1)
			 | (OP==`LDY_abs & T==`Tthree & phi2)
			 | (OP==`LDA_abs & T==`Tzero & phi1)
			 | (OP==`LDA_abs & T==`Tzero & phi2)
			 | (OP==`LDA_abs & T==`Tone & phi1)
			 | (OP==`LDA_abs & T==`Tone & phi2)
			 | (OP==`LDA_abs & T==`Ttwo & phi1)
			 | (OP==`LDA_abs & T==`Ttwo & phi2)
			 | (OP==`LDA_abs & T==`Tthree & phi1)
			 | (OP==`LDA_abs & T==`Tthree & phi2)
			 | (OP==`LDX_abs & T==`Tzero & phi1)
			 | (OP==`LDX_abs & T==`Tzero & phi2)
			 | (OP==`LDX_abs & T==`Tone & phi1)
			 | (OP==`LDX_abs & T==`Tone & phi2)
			 | (OP==`LDX_abs & T==`Ttwo & phi1)
			 | (OP==`LDX_abs & T==`Ttwo & phi2)
			 | (OP==`LDX_abs & T==`Tthree & phi1)
			 | (OP==`LDX_abs & T==`Tthree & phi2)
			 | (OP==`BCS_rel & T==`Tzero & phi1)
			 | (OP==`BCS_rel & T==`Tzero & phi2)
			 | (OP==`BCS_rel & T==`Ttwo & phi1)
			 | (OP==`BCS_rel & T==`Ttwo & phi2)
			 | (OP==`BCS_rel & T==`Tthree & phi1)
			 | (OP==`BCS_rel & T==`Tthree & phi2)
			 | (OP==`BCS_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BCS_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BCS_rel & T==`T1BranchCross & phi1)
			 | (OP==`BCS_rel & T==`T1BranchCross & phi2)
			 | (OP==`BCS_rel & T==`T1NoBranch & phi1)
			 | (OP==`BCS_rel & T==`T1NoBranch & phi2)
			 | (OP==`LDA_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDA_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`LDA_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`LDA_izy & T==`TzeroCrossPg & phi2)
			 | (OP==`LDA_izy & T==`Tone & phi1)
			 | (OP==`LDA_izy & T==`Tone & phi2)
			 | (OP==`LDA_izy & T==`Ttwo & phi1)
			 | (OP==`LDA_izy & T==`Ttwo & phi2)
			 | (OP==`LDA_izy & T==`Tthree & phi1)
			 | (OP==`LDA_izy & T==`Tthree & phi2)
			 | (OP==`LDA_izy & T==`Tfour & phi1)
			 | (OP==`LDA_izy & T==`Tfour & phi2)
			 | (OP==`LDA_izy & T==`Tfive & phi1)
			 | (OP==`LDA_izy & T==`Tfive & phi2)
			 | (OP==`LDY_zpx & T==`Tzero & phi1)
			 | (OP==`LDY_zpx & T==`Tzero & phi2)
			 | (OP==`LDY_zpx & T==`Tone & phi1)
			 | (OP==`LDY_zpx & T==`Tone & phi2)
			 | (OP==`LDY_zpx & T==`Ttwo & phi1)
			 | (OP==`LDY_zpx & T==`Ttwo & phi2)
			 | (OP==`LDY_zpx & T==`Tthree & phi1)
			 | (OP==`LDY_zpx & T==`Tthree & phi2)
			 | (OP==`LDA_zpx & T==`Tzero & phi1)
			 | (OP==`LDA_zpx & T==`Tzero & phi2)
			 | (OP==`LDA_zpx & T==`Tone & phi1)
			 | (OP==`LDA_zpx & T==`Tone & phi2)
			 | (OP==`LDA_zpx & T==`Ttwo & phi1)
			 | (OP==`LDA_zpx & T==`Ttwo & phi2)
			 | (OP==`LDA_zpx & T==`Tthree & phi1)
			 | (OP==`LDA_zpx & T==`Tthree & phi2)
			 | (OP==`LDX_zpy & T==`Tzero & phi1)
			 | (OP==`LDX_zpy & T==`Tzero & phi2)
			 | (OP==`LDX_zpy & T==`Tone & phi1)
			 | (OP==`LDX_zpy & T==`Tone & phi2)
			 | (OP==`LDX_zpy & T==`Ttwo & phi1)
			 | (OP==`LDX_zpy & T==`Ttwo & phi2)
			 | (OP==`LDX_zpy & T==`Tthree & phi1)
			 | (OP==`LDX_zpy & T==`Tthree & phi2)
			 | (OP==`CLV & T==`Tone & phi1)
			 | (OP==`CLV & T==`Tone & phi2)
			 | (OP==`CLV & T==`Ttwo & phi1)
			 | (OP==`CLV & T==`Ttwo & phi2)
			 | (OP==`LDA_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDA_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`LDA_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`LDA_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`LDA_aby & T==`Tone & phi1)
			 | (OP==`LDA_aby & T==`Tone & phi2)
			 | (OP==`LDA_aby & T==`Ttwo & phi1)
			 | (OP==`LDA_aby & T==`Ttwo & phi2)
			 | (OP==`LDA_aby & T==`Tthree & phi1)
			 | (OP==`LDA_aby & T==`Tthree & phi2)
			 | (OP==`LDA_aby & T==`Tfour & phi1)
			 | (OP==`LDA_aby & T==`Tfour & phi2)
			 | (OP==`TSX & T==`Tone & phi1)
			 | (OP==`TSX & T==`Tone & phi2)
			 | (OP==`TSX & T==`Ttwo & phi1)
			 | (OP==`TSX & T==`Ttwo & phi2)
			 | (OP==`LDY_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDY_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`LDY_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`LDY_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`LDY_abx & T==`Tone & phi1)
			 | (OP==`LDY_abx & T==`Tone & phi2)
			 | (OP==`LDY_abx & T==`Ttwo & phi1)
			 | (OP==`LDY_abx & T==`Ttwo & phi2)
			 | (OP==`LDY_abx & T==`Tthree & phi1)
			 | (OP==`LDY_abx & T==`Tthree & phi2)
			 | (OP==`LDY_abx & T==`Tfour & phi1)
			 | (OP==`LDY_abx & T==`Tfour & phi2)
			 | (OP==`LDA_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDA_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`LDA_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`LDA_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`LDA_abx & T==`Tone & phi1)
			 | (OP==`LDA_abx & T==`Tone & phi2)
			 | (OP==`LDA_abx & T==`Ttwo & phi1)
			 | (OP==`LDA_abx & T==`Ttwo & phi2)
			 | (OP==`LDA_abx & T==`Tthree & phi1)
			 | (OP==`LDA_abx & T==`Tthree & phi2)
			 | (OP==`LDA_abx & T==`Tfour & phi1)
			 | (OP==`LDA_abx & T==`Tfour & phi2)
			 | (OP==`LDX_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDX_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`LDX_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`LDX_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`LDX_aby & T==`Tone & phi1)
			 | (OP==`LDX_aby & T==`Tone & phi2)
			 | (OP==`LDX_aby & T==`Ttwo & phi1)
			 | (OP==`LDX_aby & T==`Ttwo & phi2)
			 | (OP==`LDX_aby & T==`Tthree & phi1)
			 | (OP==`LDX_aby & T==`Tthree & phi2)
			 | (OP==`LDX_aby & T==`Tfour & phi1)
			 | (OP==`LDX_aby & T==`Tfour & phi2)
			 | (OP==`CPY_imm & T==`Tone & phi1)
			 | (OP==`CPY_imm & T==`Tone & phi2)
			 | (OP==`CPY_imm & T==`Ttwo & phi1)
			 | (OP==`CPY_imm & T==`Ttwo & phi2)
			 | (OP==`CMP_izx & T==`Tzero & phi1)
			 | (OP==`CMP_izx & T==`Tzero & phi2)
			 | (OP==`CMP_izx & T==`Tone & phi1)
			 | (OP==`CMP_izx & T==`Tone & phi2)
			 | (OP==`CMP_izx & T==`Ttwo & phi1)
			 | (OP==`CMP_izx & T==`Ttwo & phi2)
			 | (OP==`CMP_izx & T==`Tthree & phi1)
			 | (OP==`CMP_izx & T==`Tthree & phi2)
			 | (OP==`CMP_izx & T==`Tfour & phi1)
			 | (OP==`CMP_izx & T==`Tfour & phi2)
			 | (OP==`CMP_izx & T==`Tfive & phi1)
			 | (OP==`CMP_izx & T==`Tfive & phi2)
			 | (OP==`CPY_zp & T==`Tzero & phi1)
			 | (OP==`CPY_zp & T==`Tzero & phi2)
			 | (OP==`CPY_zp & T==`Tone & phi1)
			 | (OP==`CPY_zp & T==`Tone & phi2)
			 | (OP==`CPY_zp & T==`Ttwo & phi1)
			 | (OP==`CPY_zp & T==`Ttwo & phi2)
			 | (OP==`CMP_zp & T==`Tzero & phi1)
			 | (OP==`CMP_zp & T==`Tzero & phi2)
			 | (OP==`CMP_zp & T==`Tone & phi1)
			 | (OP==`CMP_zp & T==`Tone & phi2)
			 | (OP==`CMP_zp & T==`Ttwo & phi1)
			 | (OP==`CMP_zp & T==`Ttwo & phi2)
			 | (OP==`DEC_zp & T==`Tzero & phi1)
			 | (OP==`DEC_zp & T==`Tzero & phi2)
			 | (OP==`DEC_zp & T==`Tone & phi1)
			 | (OP==`DEC_zp & T==`Tone & phi2)
			 | (OP==`DEC_zp & T==`Ttwo & phi1)
			 | (OP==`DEC_zp & T==`Ttwo & phi2)
			 | (OP==`DEC_zp & T==`Tthree & phi1)
			 | (OP==`DEC_zp & T==`Tthree & phi2)
			 | (OP==`DEC_zp & T==`Tfour & phi1)
			 | (OP==`DEC_zp & T==`Tfour & phi2)
			 | (OP==`INY & T==`Tone & phi1)
			 | (OP==`INY & T==`Tone & phi2)
			 | (OP==`INY & T==`Ttwo & phi1)
			 | (OP==`INY & T==`Ttwo & phi2)
			 | (OP==`CMP_imm & T==`Tone & phi1)
			 | (OP==`CMP_imm & T==`Tone & phi2)
			 | (OP==`CMP_imm & T==`Ttwo & phi1)
			 | (OP==`CMP_imm & T==`Ttwo & phi2)
			 | (OP==`DEX & T==`Tone & phi1)
			 | (OP==`DEX & T==`Tone & phi2)
			 | (OP==`DEX & T==`Ttwo & phi1)
			 | (OP==`DEX & T==`Ttwo & phi2)
			 | (OP==`CPY_abs & T==`Tzero & phi1)
			 | (OP==`CPY_abs & T==`Tzero & phi2)
			 | (OP==`CPY_abs & T==`Tone & phi1)
			 | (OP==`CPY_abs & T==`Tone & phi2)
			 | (OP==`CPY_abs & T==`Ttwo & phi1)
			 | (OP==`CPY_abs & T==`Ttwo & phi2)
			 | (OP==`CPY_abs & T==`Tthree & phi1)
			 | (OP==`CPY_abs & T==`Tthree & phi2)
			 | (OP==`CMP_abs & T==`Tzero & phi1)
			 | (OP==`CMP_abs & T==`Tzero & phi2)
			 | (OP==`CMP_abs & T==`Tone & phi1)
			 | (OP==`CMP_abs & T==`Tone & phi2)
			 | (OP==`CMP_abs & T==`Ttwo & phi1)
			 | (OP==`CMP_abs & T==`Ttwo & phi2)
			 | (OP==`CMP_abs & T==`Tthree & phi1)
			 | (OP==`CMP_abs & T==`Tthree & phi2)
			 | (OP==`DEC_abs & T==`Tzero & phi1)
			 | (OP==`DEC_abs & T==`Tzero & phi2)
			 | (OP==`DEC_abs & T==`Tone & phi1)
			 | (OP==`DEC_abs & T==`Tone & phi2)
			 | (OP==`DEC_abs & T==`Ttwo & phi1)
			 | (OP==`DEC_abs & T==`Ttwo & phi2)
			 | (OP==`DEC_abs & T==`Tthree & phi1)
			 | (OP==`DEC_abs & T==`Tthree & phi2)
			 | (OP==`DEC_abs & T==`Tfour & phi1)
			 | (OP==`DEC_abs & T==`Tfour & phi2)
			 | (OP==`DEC_abs & T==`Tfive & phi1)
			 | (OP==`DEC_abs & T==`Tfive & phi2)
			 | (OP==`BNE_rel & T==`Tzero & phi1)
			 | (OP==`BNE_rel & T==`Tzero & phi2)
			 | (OP==`BNE_rel & T==`Ttwo & phi1)
			 | (OP==`BNE_rel & T==`Ttwo & phi2)
			 | (OP==`BNE_rel & T==`Tthree & phi1)
			 | (OP==`BNE_rel & T==`Tthree & phi2)
			 | (OP==`BNE_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BNE_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BNE_rel & T==`T1BranchCross & phi1)
			 | (OP==`BNE_rel & T==`T1BranchCross & phi2)
			 | (OP==`BNE_rel & T==`T1NoBranch & phi1)
			 | (OP==`BNE_rel & T==`T1NoBranch & phi2)
			 | (OP==`CMP_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`CMP_izy & T==`TzeroCrossPg & phi2)
			 | (OP==`CMP_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`CMP_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`CMP_izy & T==`Tone & phi1)
			 | (OP==`CMP_izy & T==`Tone & phi2)
			 | (OP==`CMP_izy & T==`Ttwo & phi1)
			 | (OP==`CMP_izy & T==`Ttwo & phi2)
			 | (OP==`CMP_izy & T==`Tthree & phi1)
			 | (OP==`CMP_izy & T==`Tthree & phi2)
			 | (OP==`CMP_izy & T==`Tfour & phi1)
			 | (OP==`CMP_izy & T==`Tfour & phi2)
			 | (OP==`CMP_izy & T==`Tfive & phi1)
			 | (OP==`CMP_izy & T==`Tfive & phi2)
			 | (OP==`CMP_zpx & T==`Tzero & phi1)
			 | (OP==`CMP_zpx & T==`Tzero & phi2)
			 | (OP==`CMP_zpx & T==`Tone & phi1)
			 | (OP==`CMP_zpx & T==`Tone & phi2)
			 | (OP==`CMP_zpx & T==`Ttwo & phi1)
			 | (OP==`CMP_zpx & T==`Ttwo & phi2)
			 | (OP==`CMP_zpx & T==`Tthree & phi1)
			 | (OP==`CMP_zpx & T==`Tthree & phi2)
			 | (OP==`DEC_zpx & T==`Tzero & phi1)
			 | (OP==`DEC_zpx & T==`Tzero & phi2)
			 | (OP==`DEC_zpx & T==`Tone & phi1)
			 | (OP==`DEC_zpx & T==`Tone & phi2)
			 | (OP==`DEC_zpx & T==`Ttwo & phi1)
			 | (OP==`DEC_zpx & T==`Ttwo & phi2)
			 | (OP==`DEC_zpx & T==`Tthree & phi1)
			 | (OP==`DEC_zpx & T==`Tthree & phi2)
			 | (OP==`DEC_zpx & T==`Tfour & phi1)
			 | (OP==`DEC_zpx & T==`Tfour & phi2)
			 | (OP==`DEC_zpx & T==`Tfive & phi1)
			 | (OP==`DEC_zpx & T==`Tfive & phi2)
			 | (OP==`CLD & T==`Tone & phi1)
			 | (OP==`CLD & T==`Tone & phi2)
			 | (OP==`CLD & T==`Ttwo & phi1)
			 | (OP==`CLD & T==`Ttwo & phi2)
			 | (OP==`CMP_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`CMP_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`CMP_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`CMP_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`CMP_aby & T==`Tone & phi1)
			 | (OP==`CMP_aby & T==`Tone & phi2)
			 | (OP==`CMP_aby & T==`Ttwo & phi1)
			 | (OP==`CMP_aby & T==`Ttwo & phi2)
			 | (OP==`CMP_aby & T==`Tthree & phi1)
			 | (OP==`CMP_aby & T==`Tthree & phi2)
			 | (OP==`CMP_aby & T==`Tfour & phi1)
			 | (OP==`CMP_aby & T==`Tfour & phi2)
			 | (OP==`CMP_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`CMP_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`CMP_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`CMP_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`CMP_abx & T==`Tone & phi1)
			 | (OP==`CMP_abx & T==`Tone & phi2)
			 | (OP==`CMP_abx & T==`Ttwo & phi1)
			 | (OP==`CMP_abx & T==`Ttwo & phi2)
			 | (OP==`CMP_abx & T==`Tthree & phi1)
			 | (OP==`CMP_abx & T==`Tthree & phi2)
			 | (OP==`CMP_abx & T==`Tfour & phi1)
			 | (OP==`CMP_abx & T==`Tfour & phi2)
			 | (OP==`DEC_abx & T==`Tzero & phi1)
			 | (OP==`DEC_abx & T==`Tzero & phi2)
			 | (OP==`DEC_abx & T==`Tone & phi1)
			 | (OP==`DEC_abx & T==`Tone & phi2)
			 | (OP==`DEC_abx & T==`Ttwo & phi1)
			 | (OP==`DEC_abx & T==`Ttwo & phi2)
			 | (OP==`DEC_abx & T==`Tthree & phi1)
			 | (OP==`DEC_abx & T==`Tthree & phi2)
			 | (OP==`DEC_abx & T==`Tfour & phi1)
			 | (OP==`DEC_abx & T==`Tfour & phi2)
			 | (OP==`DEC_abx & T==`Tfive & phi1)
			 | (OP==`DEC_abx & T==`Tfive & phi2)
			 | (OP==`DEC_abx & T==`Tsix & phi1)
			 | (OP==`DEC_abx & T==`Tsix & phi2)
			 | (OP==`CPX_imm & T==`Tone & phi1)
			 | (OP==`CPX_imm & T==`Tone & phi2)
			 | (OP==`CPX_imm & T==`Ttwo & phi1)
			 | (OP==`CPX_imm & T==`Ttwo & phi2)
			 | (OP==`SBC_izx & T==`Tzero & phi1)
			 | (OP==`SBC_izx & T==`Tzero & phi2)
			 | (OP==`SBC_izx & T==`Tone & phi1)
			 | (OP==`SBC_izx & T==`Tone & phi2)
			 | (OP==`SBC_izx & T==`Ttwo & phi1)
			 | (OP==`SBC_izx & T==`Ttwo & phi2)
			 | (OP==`SBC_izx & T==`Tthree & phi1)
			 | (OP==`SBC_izx & T==`Tthree & phi2)
			 | (OP==`SBC_izx & T==`Tfour & phi1)
			 | (OP==`SBC_izx & T==`Tfour & phi2)
			 | (OP==`SBC_izx & T==`Tfive & phi1)
			 | (OP==`SBC_izx & T==`Tfive & phi2)
			 | (OP==`CPX_zp & T==`Tzero & phi1)
			 | (OP==`CPX_zp & T==`Tzero & phi2)
			 | (OP==`CPX_zp & T==`Tone & phi1)
			 | (OP==`CPX_zp & T==`Tone & phi2)
			 | (OP==`CPX_zp & T==`Ttwo & phi1)
			 | (OP==`CPX_zp & T==`Ttwo & phi2)
			 | (OP==`SBC_zp & T==`Tzero & phi1)
			 | (OP==`SBC_zp & T==`Tzero & phi2)
			 | (OP==`SBC_zp & T==`Tone & phi1)
			 | (OP==`SBC_zp & T==`Tone & phi2)
			 | (OP==`SBC_zp & T==`Ttwo & phi1)
			 | (OP==`SBC_zp & T==`Ttwo & phi2)
			 | (OP==`INC_zp & T==`Tzero & phi1)
			 | (OP==`INC_zp & T==`Tzero & phi2)
			 | (OP==`INC_zp & T==`Tone & phi1)
			 | (OP==`INC_zp & T==`Tone & phi2)
			 | (OP==`INC_zp & T==`Ttwo & phi1)
			 | (OP==`INC_zp & T==`Ttwo & phi2)
			 | (OP==`INC_zp & T==`Tthree & phi1)
			 | (OP==`INC_zp & T==`Tthree & phi2)
			 | (OP==`INC_zp & T==`Tfour & phi1)
			 | (OP==`INC_zp & T==`Tfour & phi2)
			 | (OP==`INX & T==`Tone & phi1)
			 | (OP==`INX & T==`Tone & phi2)
			 | (OP==`INX & T==`Ttwo & phi1)
			 | (OP==`INX & T==`Ttwo & phi2)
			 | (OP==`SBC_imm & T==`Tone & phi1)
			 | (OP==`SBC_imm & T==`Tone & phi2)
			 | (OP==`SBC_imm & T==`Ttwo & phi1)
			 | (OP==`SBC_imm & T==`Ttwo & phi2)
			 | (OP==`NOP & T==`Tone & phi1)
			 | (OP==`NOP & T==`Tone & phi2)
			 | (OP==`NOP & T==`Ttwo & phi1)
			 | (OP==`NOP & T==`Ttwo & phi2)
			 | (OP==`CPX_abs & T==`Tzero & phi1)
			 | (OP==`CPX_abs & T==`Tzero & phi2)
			 | (OP==`CPX_abs & T==`Tone & phi1)
			 | (OP==`CPX_abs & T==`Tone & phi2)
			 | (OP==`CPX_abs & T==`Ttwo & phi1)
			 | (OP==`CPX_abs & T==`Ttwo & phi2)
			 | (OP==`CPX_abs & T==`Tthree & phi1)
			 | (OP==`CPX_abs & T==`Tthree & phi2)
			 | (OP==`SBC_abs & T==`Tzero & phi1)
			 | (OP==`SBC_abs & T==`Tzero & phi2)
			 | (OP==`SBC_abs & T==`Tone & phi1)
			 | (OP==`SBC_abs & T==`Tone & phi2)
			 | (OP==`SBC_abs & T==`Ttwo & phi1)
			 | (OP==`SBC_abs & T==`Ttwo & phi2)
			 | (OP==`SBC_abs & T==`Tthree & phi1)
			 | (OP==`SBC_abs & T==`Tthree & phi2)
			 | (OP==`INC_abs & T==`Tzero & phi1)
			 | (OP==`INC_abs & T==`Tzero & phi2)
			 | (OP==`INC_abs & T==`Tone & phi1)
			 | (OP==`INC_abs & T==`Tone & phi2)
			 | (OP==`INC_abs & T==`Ttwo & phi1)
			 | (OP==`INC_abs & T==`Ttwo & phi2)
			 | (OP==`INC_abs & T==`Tthree & phi1)
			 | (OP==`INC_abs & T==`Tthree & phi2)
			 | (OP==`INC_abs & T==`Tfour & phi1)
			 | (OP==`INC_abs & T==`Tfour & phi2)
			 | (OP==`INC_abs & T==`Tfive & phi1)
			 | (OP==`INC_abs & T==`Tfive & phi2)
			 | (OP==`BEQ_rel & T==`Tzero & phi1)
			 | (OP==`BEQ_rel & T==`Tzero & phi2)
			 | (OP==`BEQ_rel & T==`Ttwo & phi1)
			 | (OP==`BEQ_rel & T==`Ttwo & phi2)
			 | (OP==`BEQ_rel & T==`Tthree & phi1)
			 | (OP==`BEQ_rel & T==`Tthree & phi2)
			 | (OP==`BEQ_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BEQ_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BEQ_rel & T==`T1BranchCross & phi1)
			 | (OP==`BEQ_rel & T==`T1BranchCross & phi2)
			 | (OP==`BEQ_rel & T==`T1NoBranch & phi1)
			 | (OP==`BEQ_rel & T==`T1NoBranch & phi2)
			 | (OP==`SBC_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`SBC_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`SBC_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`SBC_izy & T==`TzeroCrossPg & phi2)
			 | (OP==`SBC_izy & T==`Tone & phi1)
			 | (OP==`SBC_izy & T==`Tone & phi2)
			 | (OP==`SBC_izy & T==`Ttwo & phi1)
			 | (OP==`SBC_izy & T==`Ttwo & phi2)
			 | (OP==`SBC_izy & T==`Tthree & phi1)
			 | (OP==`SBC_izy & T==`Tthree & phi2)
			 | (OP==`SBC_izy & T==`Tfour & phi1)
			 | (OP==`SBC_izy & T==`Tfour & phi2)
			 | (OP==`SBC_izy & T==`Tfive & phi1)
			 | (OP==`SBC_izy & T==`Tfive & phi2)
			 | (OP==`SBC_zpx & T==`Tzero & phi1)
			 | (OP==`SBC_zpx & T==`Tzero & phi2)
			 | (OP==`SBC_zpx & T==`Tone & phi1)
			 | (OP==`SBC_zpx & T==`Tone & phi2)
			 | (OP==`SBC_zpx & T==`Ttwo & phi1)
			 | (OP==`SBC_zpx & T==`Ttwo & phi2)
			 | (OP==`SBC_zpx & T==`Tthree & phi1)
			 | (OP==`SBC_zpx & T==`Tthree & phi2)
			 | (OP==`INC_zpx & T==`Tzero & phi1)
			 | (OP==`INC_zpx & T==`Tzero & phi2)
			 | (OP==`INC_zpx & T==`Tone & phi1)
			 | (OP==`INC_zpx & T==`Tone & phi2)
			 | (OP==`INC_zpx & T==`Ttwo & phi1)
			 | (OP==`INC_zpx & T==`Ttwo & phi2)
			 | (OP==`INC_zpx & T==`Tthree & phi1)
			 | (OP==`INC_zpx & T==`Tthree & phi2)
			 | (OP==`INC_zpx & T==`Tfour & phi1)
			 | (OP==`INC_zpx & T==`Tfour & phi2)
			 | (OP==`INC_zpx & T==`Tfive & phi1)
			 | (OP==`INC_zpx & T==`Tfive & phi2)
			 | (OP==`SED & T==`Tone & phi1)
			 | (OP==`SED & T==`Tone & phi2)
			 | (OP==`SED & T==`Ttwo & phi1)
			 | (OP==`SED & T==`Ttwo & phi2)
			 | (OP==`SBC_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`SBC_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`SBC_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`SBC_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`SBC_aby & T==`Tone & phi1)
			 | (OP==`SBC_aby & T==`Tone & phi2)
			 | (OP==`SBC_aby & T==`Ttwo & phi1)
			 | (OP==`SBC_aby & T==`Ttwo & phi2)
			 | (OP==`SBC_aby & T==`Tthree & phi1)
			 | (OP==`SBC_aby & T==`Tthree & phi2)
			 | (OP==`SBC_aby & T==`Tfour & phi1)
			 | (OP==`SBC_aby & T==`Tfour & phi2)
			 | (OP==`SBC_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`SBC_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`SBC_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`SBC_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`SBC_abx & T==`Tone & phi1)
			 | (OP==`SBC_abx & T==`Tone & phi2)
			 | (OP==`SBC_abx & T==`Ttwo & phi1)
			 | (OP==`SBC_abx & T==`Ttwo & phi2)
			 | (OP==`SBC_abx & T==`Tthree & phi1)
			 | (OP==`SBC_abx & T==`Tthree & phi2)
			 | (OP==`SBC_abx & T==`Tfour & phi1)
			 | (OP==`SBC_abx & T==`Tfour & phi2)
			 | (OP==`INC_abx & T==`Tzero & phi1)
			 | (OP==`INC_abx & T==`Tzero & phi2)
			 | (OP==`INC_abx & T==`Tone & phi1)
			 | (OP==`INC_abx & T==`Tone & phi2)
			 | (OP==`INC_abx & T==`Ttwo & phi1)
			 | (OP==`INC_abx & T==`Ttwo & phi2)
			 | (OP==`INC_abx & T==`Tthree & phi1)
			 | (OP==`INC_abx & T==`Tthree & phi2)
			 | (OP==`INC_abx & T==`Tfour & phi1)
			 | (OP==`INC_abx & T==`Tfour & phi2)
			 | (OP==`INC_abx & T==`Tfive & phi1)
			 | (OP==`INC_abx & T==`Tfive & phi2)
			 | (OP==`INC_abx & T==`Tsix & phi1)
			 | (OP==`INC_abx & T==`Tsix & phi2)
			;

assign control[`ANDS] = (OP==`AND_izx & T==`Tone & phi1)
			 | (OP==`AND_izx & T==`Tone & phi2)
			 | (OP==`BIT_zp & T==`Tone & phi1)
			 | (OP==`BIT_zp & T==`Tone & phi2)
			 | (OP==`AND_zp & T==`Tone & phi1)
			 | (OP==`AND_zp & T==`Tone & phi2)
			 | (OP==`AND_imm & T==`Tone & phi1)
			 | (OP==`AND_imm & T==`Tone & phi2)
			 | (OP==`BIT_abs & T==`Tone & phi1)
			 | (OP==`BIT_abs & T==`Tone & phi2)
			 | (OP==`AND_abs & T==`Tone & phi1)
			 | (OP==`AND_abs & T==`Tone & phi2)
			 | (OP==`AND_izy & T==`Tone & phi1)
			 | (OP==`AND_izy & T==`Tone & phi2)
			 | (OP==`AND_zpx & T==`Tone & phi1)
			 | (OP==`AND_zpx & T==`Tone & phi2)
			 | (OP==`AND_aby & T==`Tone & phi1)
			 | (OP==`AND_aby & T==`Tone & phi2)
			 | (OP==`AND_abx & T==`Tone & phi1)
			 | (OP==`AND_abx & T==`Tone & phi2)
			;

assign control[`EORS] = (OP==`EOR_izx & T==`Tone & phi1)
			 | (OP==`EOR_izx & T==`Tone & phi2)
			 | (OP==`EOR_zp & T==`Tone & phi1)
			 | (OP==`EOR_zp & T==`Tone & phi2)
			 | (OP==`EOR_imm & T==`Tone & phi1)
			 | (OP==`EOR_imm & T==`Tone & phi2)
			 | (OP==`EOR_abs & T==`Tone & phi1)
			 | (OP==`EOR_abs & T==`Tone & phi2)
			 | (OP==`EOR_izy & T==`Tone & phi1)
			 | (OP==`EOR_izy & T==`Tone & phi2)
			 | (OP==`EOR_zpx & T==`Tone & phi1)
			 | (OP==`EOR_zpx & T==`Tone & phi2)
			 | (OP==`EOR_aby & T==`Tone & phi1)
			 | (OP==`EOR_aby & T==`Tone & phi2)
			 | (OP==`EOR_abx & T==`Tone & phi1)
			 | (OP==`EOR_abx & T==`Tone & phi2)
			;

assign control[`ORS] = (OP==`ORA_izx & T==`Tone & phi1)
			 | (OP==`ORA_izx & T==`Tone & phi2)
			 | (OP==`ORA_zp & T==`Tone & phi1)
			 | (OP==`ORA_zp & T==`Tone & phi2)
			 | (OP==`ORA_imm & T==`Tone & phi1)
			 | (OP==`ORA_imm & T==`Tone & phi2)
			 | (OP==`ORA_abs & T==`Tone & phi1)
			 | (OP==`ORA_abs & T==`Tone & phi2)
			 | (OP==`ASL_abs & T==`Tone & phi2)
			 | (OP==`ORA_izy & T==`Tone & phi1)
			 | (OP==`ORA_izy & T==`Tone & phi2)
			 | (OP==`ORA_zpx & T==`Tone & phi1)
			 | (OP==`ORA_zpx & T==`Tone & phi2)
			 | (OP==`ORA_aby & T==`Tone & phi1)
			 | (OP==`ORA_aby & T==`Tone & phi2)
			 | (OP==`ORA_abx & T==`Tone & phi1)
			 | (OP==`ORA_abx & T==`Tone & phi2)
			;

assign control[`SRS] = (OP==`LSR_zp & T==`Tfour & phi1)
			 | (OP==`LSR_zp & T==`Tfour & phi2)
			 | (OP==`LSR & T==`Tone & phi1)
			 | (OP==`LSR & T==`Tone & phi2)
			 | (OP==`LSR_abs & T==`Tfive & phi1)
			 | (OP==`LSR_abs & T==`Tfive & phi2)
			 | (OP==`LSR_zpx & T==`Tfive & phi1)
			 | (OP==`LSR_zpx & T==`Tfive & phi2)
			 | (OP==`LSR_abx & T==`Tsix & phi1)
			 | (OP==`LSR_abx & T==`Tsix & phi2)
			 | (OP==`ROR_zp & T==`Tfour & phi1)
			 | (OP==`ROR_zp & T==`Tfour & phi2)
			 | (OP==`ROR & T==`Tone & phi1)
			 | (OP==`ROR & T==`Tone & phi2)
			 | (OP==`ROR_abs & T==`Tfive & phi1)
			 | (OP==`ROR_abs & T==`Tfive & phi2)
			 | (OP==`ROR_zpx & T==`Tfive & phi1)
			 | (OP==`ROR_zpx & T==`Tfive & phi2)
			 | (OP==`ROR_abx & T==`Tsix & phi1)
			 | (OP==`ROR_abx & T==`Tsix & phi2)
			;

assign control[`ADD_ADL] = (OP==`BRK & T==`Tzero & phi2)
			 | (OP==`BRK & T==`Tone & phi1)
			 | (OP==`BRK & T==`Tthree & phi2)
			 | (OP==`BRK & T==`Tfour & phi1)
			 | (OP==`BRK & T==`Tfour & phi2)
			 | (OP==`BRK & T==`Tfive & phi1)
			 | (OP==`ORA_izx & T==`Tzero & phi1)
			 | (OP==`ORA_izx & T==`Tthree & phi2)
			 | (OP==`ORA_izx & T==`Tfour & phi1)
			 | (OP==`ORA_izx & T==`Tfour & phi2)
			 | (OP==`ORA_izx & T==`Tfive & phi1)
			 | (OP==`ORA_izx & T==`Tfive & phi2)
			 | (OP==`ASL_zp & T==`Tzero & phi1)
			 | (OP==`ASL_zp & T==`Tthree & phi2)
			 | (OP==`ASL_zp & T==`Tfour & phi1)
			 | (OP==`ASL_zp & T==`Tfour & phi2)
			 | (OP==`ORA_abs & T==`Tzero & phi1)
			 | (OP==`ORA_abs & T==`Tthree & phi2)
			 | (OP==`ASL_abs & T==`Tthree & phi2)
			 | (OP==`ASL_abs & T==`Tfour & phi1)
			 | (OP==`ASL_abs & T==`Tfour & phi2)
			 | (OP==`ASL_abs & T==`Tfive & phi1)
			 | (OP==`BPL_rel & T==`Tzero & phi1)
			 | (OP==`BPL_rel & T==`Tthree & phi2)
			 | (OP==`BPL_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`ORA_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ORA_izy & T==`Tthree & phi2)
			 | (OP==`ORA_izy & T==`Tfour & phi1)
			 | (OP==`ORA_izy & T==`Tfour & phi2)
			 | (OP==`ORA_izy & T==`Tfive & phi1)
			 | (OP==`ORA_zpx & T==`Tzero & phi1)
			 | (OP==`ORA_zpx & T==`Tthree & phi2)
			 | (OP==`ASL_zpx & T==`Tthree & phi2)
			 | (OP==`ASL_zpx & T==`Tfour & phi1)
			 | (OP==`ASL_zpx & T==`Tfour & phi2)
			 | (OP==`ASL_zpx & T==`Tfive & phi1)
			 | (OP==`ORA_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ORA_aby & T==`Tthree & phi2)
			 | (OP==`ORA_aby & T==`Tfour & phi1)
			 | (OP==`ORA_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ORA_abx & T==`Tthree & phi2)
			 | (OP==`ORA_abx & T==`Tfour & phi1)
			 | (OP==`ASL_abx & T==`Tthree & phi2)
			 | (OP==`ASL_abx & T==`Tfour & phi1)
			 | (OP==`JSR_abs & T==`Tthree & phi2)
			 | (OP==`JSR_abs & T==`Tfour & phi1)
			 | (OP==`JSR_abs & T==`Tfour & phi2)
			 | (OP==`JSR_abs & T==`Tfive & phi1)
			 | (OP==`AND_izx & T==`Tzero & phi1)
			 | (OP==`AND_izx & T==`Tthree & phi2)
			 | (OP==`AND_izx & T==`Tfour & phi1)
			 | (OP==`AND_izx & T==`Tfour & phi2)
			 | (OP==`AND_izx & T==`Tfive & phi1)
			 | (OP==`AND_izx & T==`Tfive & phi2)
			 | (OP==`ROL_zp & T==`Tzero & phi1)
			 | (OP==`ROL_zp & T==`Tthree & phi2)
			 | (OP==`ROL_zp & T==`Tfour & phi1)
			 | (OP==`ROL_zp & T==`Tfour & phi2)
			 | (OP==`PLP & T==`Tzero & phi1)
			 | (OP==`PLP & T==`Tthree & phi2)
			 | (OP==`BIT_abs & T==`Tzero & phi1)
			 | (OP==`BIT_abs & T==`Tthree & phi2)
			 | (OP==`AND_abs & T==`Tzero & phi1)
			 | (OP==`AND_abs & T==`Tthree & phi2)
			 | (OP==`ROL_abs & T==`Tthree & phi2)
			 | (OP==`ROL_abs & T==`Tfour & phi1)
			 | (OP==`ROL_abs & T==`Tfour & phi2)
			 | (OP==`ROL_abs & T==`Tfive & phi1)
			 | (OP==`BMI_rel & T==`Tzero & phi1)
			 | (OP==`BMI_rel & T==`Tthree & phi2)
			 | (OP==`BMI_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`AND_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`AND_izy & T==`Tthree & phi2)
			 | (OP==`AND_izy & T==`Tfour & phi1)
			 | (OP==`AND_izy & T==`Tfour & phi2)
			 | (OP==`AND_izy & T==`Tfive & phi1)
			 | (OP==`AND_zpx & T==`Tzero & phi1)
			 | (OP==`AND_zpx & T==`Tthree & phi2)
			 | (OP==`ROL_zpx & T==`Tthree & phi2)
			 | (OP==`ROL_zpx & T==`Tfour & phi1)
			 | (OP==`ROL_zpx & T==`Tfour & phi2)
			 | (OP==`ROL_zpx & T==`Tfive & phi1)
			 | (OP==`AND_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`AND_aby & T==`Tthree & phi2)
			 | (OP==`AND_aby & T==`Tfour & phi1)
			 | (OP==`AND_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`AND_abx & T==`Tthree & phi2)
			 | (OP==`AND_abx & T==`Tfour & phi1)
			 | (OP==`ROL_abx & T==`Tthree & phi2)
			 | (OP==`ROL_abx & T==`Tfour & phi1)
			 | (OP==`RTI & T==`Tzero & phi1)
			 | (OP==`RTI & T==`Tzero & phi2)
			 | (OP==`RTI & T==`Tone & phi1)
			 | (OP==`RTI & T==`Tthree & phi2)
			 | (OP==`RTI & T==`Tfour & phi1)
			 | (OP==`RTI & T==`Tfour & phi2)
			 | (OP==`RTI & T==`Tfive & phi1)
			 | (OP==`RTI & T==`Tfive & phi2)
			 | (OP==`EOR_izx & T==`Tzero & phi1)
			 | (OP==`EOR_izx & T==`Tthree & phi2)
			 | (OP==`EOR_izx & T==`Tfour & phi1)
			 | (OP==`EOR_izx & T==`Tfour & phi2)
			 | (OP==`EOR_izx & T==`Tfive & phi1)
			 | (OP==`EOR_izx & T==`Tfive & phi2)
			 | (OP==`LSR_zp & T==`Tzero & phi1)
			 | (OP==`LSR_zp & T==`Tthree & phi2)
			 | (OP==`LSR_zp & T==`Tfour & phi1)
			 | (OP==`LSR_zp & T==`Tfour & phi2)
			 | (OP==`JMP_abs & T==`Tzero & phi2)
			 | (OP==`JMP_abs & T==`Tone & phi1)
			 | (OP==`EOR_abs & T==`Tzero & phi1)
			 | (OP==`EOR_abs & T==`Tthree & phi2)
			 | (OP==`LSR_abs & T==`Tthree & phi2)
			 | (OP==`LSR_abs & T==`Tfour & phi1)
			 | (OP==`LSR_abs & T==`Tfour & phi2)
			 | (OP==`LSR_abs & T==`Tfive & phi1)
			 | (OP==`BVC_rel & T==`Tzero & phi1)
			 | (OP==`BVC_rel & T==`Tthree & phi2)
			 | (OP==`BVC_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`EOR_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`EOR_izy & T==`Tthree & phi2)
			 | (OP==`EOR_izy & T==`Tfour & phi1)
			 | (OP==`EOR_izy & T==`Tfour & phi2)
			 | (OP==`EOR_izy & T==`Tfive & phi1)
			 | (OP==`EOR_zpx & T==`Tzero & phi1)
			 | (OP==`EOR_zpx & T==`Tthree & phi2)
			 | (OP==`LSR_zpx & T==`Tthree & phi2)
			 | (OP==`LSR_zpx & T==`Tfour & phi1)
			 | (OP==`LSR_zpx & T==`Tfour & phi2)
			 | (OP==`LSR_zpx & T==`Tfive & phi1)
			 | (OP==`EOR_aby & T==`Tthree & phi2)
			 | (OP==`EOR_aby & T==`Tfour & phi1)
			 | (OP==`EOR_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`EOR_abx & T==`Tthree & phi2)
			 | (OP==`EOR_abx & T==`Tfour & phi1)
			 | (OP==`LSR_abx & T==`Tthree & phi2)
			 | (OP==`LSR_abx & T==`Tfour & phi1)
			 | (OP==`RTS & T==`Tzero & phi1)
			 | (OP==`RTS & T==`Tthree & phi2)
			 | (OP==`RTS & T==`Tfour & phi1)
			 | (OP==`RTS & T==`Tfour & phi2)
			 | (OP==`RTS & T==`Tfive & phi1)
			 | (OP==`RTS & T==`Tfive & phi2)
			 | (OP==`ADC_izx & T==`Tzero & phi1)
			 | (OP==`ADC_izx & T==`Tthree & phi2)
			 | (OP==`ADC_izx & T==`Tfour & phi1)
			 | (OP==`ADC_izx & T==`Tfour & phi2)
			 | (OP==`ADC_izx & T==`Tfive & phi1)
			 | (OP==`ADC_izx & T==`Tfive & phi2)
			 | (OP==`ROR_zp & T==`Tzero & phi1)
			 | (OP==`ROR_zp & T==`Tthree & phi2)
			 | (OP==`ROR_zp & T==`Tfour & phi1)
			 | (OP==`ROR_zp & T==`Tfour & phi2)
			 | (OP==`PLA & T==`Tzero & phi1)
			 | (OP==`PLA & T==`Tthree & phi2)
			 | (OP==`JMP_zp & T==`Tzero & phi1)
			 | (OP==`JMP_zp & T==`Tzero & phi2)
			 | (OP==`JMP_zp & T==`Tone & phi1)
			 | (OP==`JMP_zp & T==`Tthree & phi2)
			 | (OP==`JMP_zp & T==`Tfour & phi1)
			 | (OP==`JMP_zp & T==`Tfour & phi2)
			 | (OP==`ADC_abs & T==`Tzero & phi1)
			 | (OP==`ADC_abs & T==`Tthree & phi2)
			 | (OP==`ROR_abs & T==`Tthree & phi2)
			 | (OP==`ROR_abs & T==`Tfour & phi1)
			 | (OP==`ROR_abs & T==`Tfour & phi2)
			 | (OP==`ROR_abs & T==`Tfive & phi1)
			 | (OP==`BVS_rel & T==`Tzero & phi1)
			 | (OP==`BVS_rel & T==`Tthree & phi2)
			 | (OP==`BVS_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`ADC_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ADC_izy & T==`Tthree & phi2)
			 | (OP==`ADC_izy & T==`Tfour & phi1)
			 | (OP==`ADC_izy & T==`Tfour & phi2)
			 | (OP==`ADC_izy & T==`Tfive & phi1)
			 | (OP==`ADC_zpx & T==`Tzero & phi1)
			 | (OP==`ADC_zpx & T==`Tthree & phi2)
			 | (OP==`ROR_zpx & T==`Tthree & phi2)
			 | (OP==`ROR_zpx & T==`Tfour & phi1)
			 | (OP==`ROR_zpx & T==`Tfour & phi2)
			 | (OP==`ROR_zpx & T==`Tfive & phi1)
			 | (OP==`ADC_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ADC_aby & T==`Tthree & phi2)
			 | (OP==`ADC_aby & T==`Tfour & phi1)
			 | (OP==`ADC_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ADC_abx & T==`Tthree & phi2)
			 | (OP==`ADC_abx & T==`Tfour & phi1)
			 | (OP==`ROR_abx & T==`Tthree & phi2)
			 | (OP==`ROR_abx & T==`Tfour & phi1)
			 | (OP==`STA_izx & T==`Tzero & phi1)
			 | (OP==`STA_izx & T==`Tthree & phi2)
			 | (OP==`STA_izx & T==`Tfour & phi1)
			 | (OP==`STA_izx & T==`Tfour & phi2)
			 | (OP==`STA_izx & T==`Tfive & phi1)
			 | (OP==`STA_izx & T==`Tfive & phi2)
			 | (OP==`STY_abs & T==`Tzero & phi1)
			 | (OP==`STY_abs & T==`Tthree & phi2)
			 | (OP==`STA_abs & T==`Tzero & phi1)
			 | (OP==`STA_abs & T==`Tthree & phi2)
			 | (OP==`STX_abs & T==`Tzero & phi1)
			 | (OP==`STX_abs & T==`Tthree & phi2)
			 | (OP==`BCC_rel & T==`Tzero & phi1)
			 | (OP==`BCC_rel & T==`Tthree & phi2)
			 | (OP==`BCC_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`STA_izy & T==`Tthree & phi2)
			 | (OP==`STA_izy & T==`Tfour & phi1)
			 | (OP==`STA_izy & T==`Tfour & phi2)
			 | (OP==`STA_izy & T==`Tfive & phi1)
			 | (OP==`STY_zpx & T==`Tzero & phi1)
			 | (OP==`STY_zpx & T==`Tthree & phi2)
			 | (OP==`STA_zpx & T==`Tzero & phi1)
			 | (OP==`STA_zpx & T==`Tthree & phi2)
			 | (OP==`STX_zpy & T==`Tzero & phi1)
			 | (OP==`STX_zpy & T==`Tthree & phi2)
			 | (OP==`STA_aby & T==`Tthree & phi2)
			 | (OP==`STA_aby & T==`Tfour & phi1)
			 | (OP==`STA_abx & T==`Tthree & phi2)
			 | (OP==`STA_abx & T==`Tfour & phi1)
			 | (OP==`LDA_izx & T==`Tzero & phi1)
			 | (OP==`LDA_izx & T==`Tthree & phi2)
			 | (OP==`LDA_izx & T==`Tfour & phi1)
			 | (OP==`LDA_izx & T==`Tfour & phi2)
			 | (OP==`LDA_izx & T==`Tfive & phi1)
			 | (OP==`LDA_izx & T==`Tfive & phi2)
			 | (OP==`LDY_abs & T==`Tzero & phi1)
			 | (OP==`LDY_abs & T==`Tthree & phi2)
			 | (OP==`LDA_abs & T==`Tzero & phi1)
			 | (OP==`LDA_abs & T==`Tthree & phi2)
			 | (OP==`LDX_abs & T==`Tzero & phi1)
			 | (OP==`LDX_abs & T==`Tthree & phi2)
			 | (OP==`BCS_rel & T==`Tzero & phi1)
			 | (OP==`BCS_rel & T==`Tthree & phi2)
			 | (OP==`BCS_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`LDA_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDA_izy & T==`Tthree & phi2)
			 | (OP==`LDA_izy & T==`Tfour & phi1)
			 | (OP==`LDA_izy & T==`Tfour & phi2)
			 | (OP==`LDA_izy & T==`Tfive & phi1)
			 | (OP==`LDY_zpx & T==`Tzero & phi1)
			 | (OP==`LDY_zpx & T==`Tthree & phi2)
			 | (OP==`LDA_zpx & T==`Tzero & phi1)
			 | (OP==`LDA_zpx & T==`Tthree & phi2)
			 | (OP==`LDX_zpy & T==`Tzero & phi1)
			 | (OP==`LDX_zpy & T==`Tthree & phi2)
			 | (OP==`LDA_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDA_aby & T==`Tthree & phi2)
			 | (OP==`LDA_aby & T==`Tfour & phi1)
			 | (OP==`LDY_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDY_abx & T==`Tthree & phi2)
			 | (OP==`LDY_abx & T==`Tfour & phi1)
			 | (OP==`LDA_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDA_abx & T==`Tthree & phi2)
			 | (OP==`LDA_abx & T==`Tfour & phi1)
			 | (OP==`LDX_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDX_aby & T==`Tthree & phi2)
			 | (OP==`LDX_aby & T==`Tfour & phi1)
			 | (OP==`CMP_izx & T==`Tzero & phi1)
			 | (OP==`CMP_izx & T==`Tthree & phi2)
			 | (OP==`CMP_izx & T==`Tfour & phi1)
			 | (OP==`CMP_izx & T==`Tfour & phi2)
			 | (OP==`CMP_izx & T==`Tfive & phi1)
			 | (OP==`CMP_izx & T==`Tfive & phi2)
			 | (OP==`DEC_zp & T==`Tzero & phi1)
			 | (OP==`DEC_zp & T==`Tthree & phi2)
			 | (OP==`DEC_zp & T==`Tfour & phi1)
			 | (OP==`DEC_zp & T==`Tfour & phi2)
			 | (OP==`CPY_abs & T==`Tzero & phi1)
			 | (OP==`CPY_abs & T==`Tthree & phi2)
			 | (OP==`CMP_abs & T==`Tzero & phi1)
			 | (OP==`CMP_abs & T==`Tthree & phi2)
			 | (OP==`DEC_abs & T==`Tthree & phi2)
			 | (OP==`DEC_abs & T==`Tfour & phi1)
			 | (OP==`DEC_abs & T==`Tfour & phi2)
			 | (OP==`DEC_abs & T==`Tfive & phi1)
			 | (OP==`BNE_rel & T==`Tzero & phi1)
			 | (OP==`BNE_rel & T==`Tthree & phi2)
			 | (OP==`BNE_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`CMP_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`CMP_izy & T==`Tthree & phi2)
			 | (OP==`CMP_izy & T==`Tfour & phi1)
			 | (OP==`CMP_izy & T==`Tfour & phi2)
			 | (OP==`CMP_izy & T==`Tfive & phi1)
			 | (OP==`CMP_zpx & T==`Tzero & phi1)
			 | (OP==`CMP_zpx & T==`Tthree & phi2)
			 | (OP==`DEC_zpx & T==`Tthree & phi2)
			 | (OP==`DEC_zpx & T==`Tfour & phi1)
			 | (OP==`DEC_zpx & T==`Tfour & phi2)
			 | (OP==`DEC_zpx & T==`Tfive & phi1)
			 | (OP==`CMP_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`CMP_aby & T==`Tthree & phi2)
			 | (OP==`CMP_aby & T==`Tfour & phi1)
			 | (OP==`CMP_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`CMP_abx & T==`Tthree & phi2)
			 | (OP==`CMP_abx & T==`Tfour & phi1)
			 | (OP==`DEC_abx & T==`Tthree & phi2)
			 | (OP==`DEC_abx & T==`Tfour & phi1)
			 | (OP==`SBC_izx & T==`Tzero & phi1)
			 | (OP==`SBC_izx & T==`Tthree & phi2)
			 | (OP==`SBC_izx & T==`Tfour & phi1)
			 | (OP==`SBC_izx & T==`Tfour & phi2)
			 | (OP==`SBC_izx & T==`Tfive & phi1)
			 | (OP==`SBC_izx & T==`Tfive & phi2)
			 | (OP==`INC_zp & T==`Tzero & phi1)
			 | (OP==`INC_zp & T==`Tthree & phi2)
			 | (OP==`INC_zp & T==`Tfour & phi1)
			 | (OP==`INC_zp & T==`Tfour & phi2)
			 | (OP==`CPX_abs & T==`Tzero & phi1)
			 | (OP==`CPX_abs & T==`Tthree & phi2)
			 | (OP==`SBC_abs & T==`Tzero & phi1)
			 | (OP==`SBC_abs & T==`Tthree & phi2)
			 | (OP==`INC_abs & T==`Tthree & phi2)
			 | (OP==`INC_abs & T==`Tfour & phi1)
			 | (OP==`INC_abs & T==`Tfour & phi2)
			 | (OP==`INC_abs & T==`Tfive & phi1)
			 | (OP==`BEQ_rel & T==`Tzero & phi1)
			 | (OP==`BEQ_rel & T==`Tthree & phi2)
			 | (OP==`BEQ_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`SBC_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`SBC_izy & T==`Tthree & phi2)
			 | (OP==`SBC_izy & T==`Tfour & phi1)
			 | (OP==`SBC_izy & T==`Tfour & phi2)
			 | (OP==`SBC_izy & T==`Tfive & phi1)
			 | (OP==`SBC_zpx & T==`Tzero & phi1)
			 | (OP==`SBC_zpx & T==`Tthree & phi2)
			 | (OP==`INC_zpx & T==`Tthree & phi2)
			 | (OP==`INC_zpx & T==`Tfour & phi1)
			 | (OP==`INC_zpx & T==`Tfour & phi2)
			 | (OP==`INC_zpx & T==`Tfive & phi1)
			 | (OP==`SBC_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`SBC_aby & T==`Tthree & phi2)
			 | (OP==`SBC_aby & T==`Tfour & phi1)
			 | (OP==`SBC_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`SBC_abx & T==`Tthree & phi2)
			 | (OP==`SBC_abx & T==`Tfour & phi1)
			 | (OP==`INC_abx & T==`Tthree & phi2)
			 | (OP==`INC_abx & T==`Tfour & phi1)
			;

assign control[`ADD_SB0to6] = (OP==`BRK & T==`Tone & phi2)
			 | (OP==`BRK & T==`Ttwo & phi1)
			 | (OP==`BRK & T==`Tfive & phi2)
			 | (OP==`BRK & T==`Tsix & phi1)
			 | (OP==`ORA_izx & T==`Tone & phi2)
			 | (OP==`ORA_izx & T==`Ttwo & phi1)
			 | (OP==`ORA_zp & T==`Tone & phi2)
			 | (OP==`ORA_zp & T==`Ttwo & phi1)
			 | (OP==`ASL_zp & T==`Tzero & phi1)
			 | (OP==`ASL_zp & T==`Tone & phi2)
			 | (OP==`ASL_zp & T==`Ttwo & phi1)
			 | (OP==`ASL_zp & T==`Tfour & phi2)
			 | (OP==`PHP & T==`Tzero & phi2)
			 | (OP==`PHP & T==`Tone & phi1)
			 | (OP==`PHP & T==`Tone & phi2)
			 | (OP==`PHP & T==`Ttwo & phi1)
			 | (OP==`ORA_imm & T==`Tone & phi2)
			 | (OP==`ORA_imm & T==`Ttwo & phi1)
			 | (OP==`ASL & T==`Tone & phi2)
			 | (OP==`ASL & T==`Ttwo & phi1)
			 | (OP==`ORA_abs & T==`Tone & phi2)
			 | (OP==`ORA_abs & T==`Ttwo & phi1)
			 | (OP==`ASL_abs & T==`Tzero & phi1)
			 | (OP==`ASL_abs & T==`Tone & phi2)
			 | (OP==`ASL_abs & T==`Ttwo & phi1)
			 | (OP==`ASL_abs & T==`Tfive & phi2)
			 | (OP==`BPL_rel & T==`Tzero & phi2)
			 | (OP==`BPL_rel & T==`Ttwo & phi1)
			 | (OP==`BPL_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BPL_rel & T==`T1BranchCross & phi1)
			 | (OP==`BPL_rel & T==`T1BranchCross & phi2)
			 | (OP==`BPL_rel & T==`T1NoBranch & phi2)
			 | (OP==`ORA_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`ORA_izy & T==`Tone & phi2)
			 | (OP==`ORA_izy & T==`Ttwo & phi1)
			 | (OP==`ORA_izy & T==`Tfive & phi2)
			 | (OP==`ORA_zpx & T==`Tone & phi2)
			 | (OP==`ORA_zpx & T==`Ttwo & phi1)
			 | (OP==`ASL_zpx & T==`Tzero & phi1)
			 | (OP==`ASL_zpx & T==`Tone & phi2)
			 | (OP==`ASL_zpx & T==`Ttwo & phi1)
			 | (OP==`ASL_zpx & T==`Tfive & phi2)
			 | (OP==`CLC & T==`Tone & phi2)
			 | (OP==`CLC & T==`Ttwo & phi1)
			 | (OP==`ORA_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`ORA_aby & T==`Tone & phi2)
			 | (OP==`ORA_aby & T==`Ttwo & phi1)
			 | (OP==`ORA_aby & T==`Tfour & phi2)
			 | (OP==`ORA_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`ORA_abx & T==`Tone & phi2)
			 | (OP==`ORA_abx & T==`Ttwo & phi1)
			 | (OP==`ORA_abx & T==`Tfour & phi2)
			 | (OP==`ASL_abx & T==`Tzero & phi1)
			 | (OP==`ASL_abx & T==`Tone & phi2)
			 | (OP==`ASL_abx & T==`Ttwo & phi1)
			 | (OP==`ASL_abx & T==`Tfour & phi2)
			 | (OP==`ASL_abx & T==`Tfive & phi1)
			 | (OP==`ASL_abx & T==`Tsix & phi2)
			 | (OP==`JSR_abs & T==`Tzero & phi1)
			 | (OP==`JSR_abs & T==`Tzero & phi2)
			 | (OP==`JSR_abs & T==`Tone & phi1)
			 | (OP==`JSR_abs & T==`Tone & phi2)
			 | (OP==`JSR_abs & T==`Ttwo & phi1)
			 | (OP==`JSR_abs & T==`Tfive & phi2)
			 | (OP==`AND_izx & T==`Tone & phi2)
			 | (OP==`AND_izx & T==`Ttwo & phi1)
			 | (OP==`BIT_zp & T==`Tone & phi2)
			 | (OP==`BIT_zp & T==`Ttwo & phi1)
			 | (OP==`AND_zp & T==`Tone & phi2)
			 | (OP==`AND_zp & T==`Ttwo & phi1)
			 | (OP==`ROL_zp & T==`Tzero & phi1)
			 | (OP==`ROL_zp & T==`Tone & phi2)
			 | (OP==`ROL_zp & T==`Ttwo & phi1)
			 | (OP==`ROL_zp & T==`Tfour & phi2)
			 | (OP==`PLP & T==`Tzero & phi1)
			 | (OP==`PLP & T==`Tone & phi2)
			 | (OP==`PLP & T==`Ttwo & phi1)
			 | (OP==`PLP & T==`Tthree & phi2)
			 | (OP==`AND_imm & T==`Tone & phi2)
			 | (OP==`AND_imm & T==`Ttwo & phi1)
			 | (OP==`ROL & T==`Tone & phi2)
			 | (OP==`ROL & T==`Ttwo & phi1)
			 | (OP==`BIT_abs & T==`Tone & phi2)
			 | (OP==`BIT_abs & T==`Ttwo & phi1)
			 | (OP==`AND_abs & T==`Tone & phi2)
			 | (OP==`AND_abs & T==`Ttwo & phi1)
			 | (OP==`ROL_abs & T==`Tzero & phi1)
			 | (OP==`ROL_abs & T==`Tone & phi2)
			 | (OP==`ROL_abs & T==`Ttwo & phi1)
			 | (OP==`ROL_abs & T==`Tfive & phi2)
			 | (OP==`BMI_rel & T==`Tzero & phi2)
			 | (OP==`BMI_rel & T==`Ttwo & phi1)
			 | (OP==`BMI_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BMI_rel & T==`T1BranchCross & phi1)
			 | (OP==`BMI_rel & T==`T1BranchCross & phi2)
			 | (OP==`BMI_rel & T==`T1NoBranch & phi2)
			 | (OP==`AND_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`AND_izy & T==`Tone & phi2)
			 | (OP==`AND_izy & T==`Ttwo & phi1)
			 | (OP==`AND_izy & T==`Tfive & phi2)
			 | (OP==`AND_zpx & T==`Tone & phi2)
			 | (OP==`AND_zpx & T==`Ttwo & phi1)
			 | (OP==`ROL_zpx & T==`Tzero & phi1)
			 | (OP==`ROL_zpx & T==`Tone & phi2)
			 | (OP==`ROL_zpx & T==`Ttwo & phi1)
			 | (OP==`ROL_zpx & T==`Tfive & phi2)
			 | (OP==`SEC & T==`Tone & phi2)
			 | (OP==`SEC & T==`Ttwo & phi1)
			 | (OP==`AND_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`AND_aby & T==`Tone & phi2)
			 | (OP==`AND_aby & T==`Ttwo & phi1)
			 | (OP==`AND_aby & T==`Tfour & phi2)
			 | (OP==`AND_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`AND_abx & T==`Tone & phi2)
			 | (OP==`AND_abx & T==`Ttwo & phi1)
			 | (OP==`AND_abx & T==`Tfour & phi2)
			 | (OP==`ROL_abx & T==`Tzero & phi1)
			 | (OP==`ROL_abx & T==`Tone & phi2)
			 | (OP==`ROL_abx & T==`Ttwo & phi1)
			 | (OP==`ROL_abx & T==`Tfour & phi2)
			 | (OP==`ROL_abx & T==`Tfive & phi1)
			 | (OP==`ROL_abx & T==`Tsix & phi2)
			 | (OP==`RTI & T==`Tzero & phi1)
			 | (OP==`RTI & T==`Tone & phi2)
			 | (OP==`RTI & T==`Ttwo & phi1)
			 | (OP==`RTI & T==`Tfive & phi2)
			 | (OP==`EOR_izx & T==`Tone & phi2)
			 | (OP==`EOR_izx & T==`Ttwo & phi1)
			 | (OP==`EOR_zp & T==`Tone & phi2)
			 | (OP==`EOR_zp & T==`Ttwo & phi1)
			 | (OP==`LSR_zp & T==`Tzero & phi1)
			 | (OP==`LSR_zp & T==`Tone & phi2)
			 | (OP==`LSR_zp & T==`Ttwo & phi1)
			 | (OP==`LSR_zp & T==`Tfour & phi2)
			 | (OP==`PHA & T==`Tzero & phi2)
			 | (OP==`PHA & T==`Tone & phi1)
			 | (OP==`PHA & T==`Tone & phi2)
			 | (OP==`PHA & T==`Ttwo & phi1)
			 | (OP==`EOR_imm & T==`Tone & phi2)
			 | (OP==`EOR_imm & T==`Ttwo & phi1)
			 | (OP==`LSR & T==`Tone & phi2)
			 | (OP==`LSR & T==`Ttwo & phi1)
			 | (OP==`JMP_abs & T==`Tone & phi2)
			 | (OP==`JMP_abs & T==`Ttwo & phi1)
			 | (OP==`EOR_abs & T==`Tone & phi2)
			 | (OP==`EOR_abs & T==`Ttwo & phi1)
			 | (OP==`LSR_abs & T==`Tzero & phi1)
			 | (OP==`LSR_abs & T==`Tone & phi2)
			 | (OP==`LSR_abs & T==`Ttwo & phi1)
			 | (OP==`LSR_abs & T==`Tfive & phi2)
			 | (OP==`BVC_rel & T==`Tzero & phi2)
			 | (OP==`BVC_rel & T==`Ttwo & phi1)
			 | (OP==`BVC_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BVC_rel & T==`T1BranchCross & phi1)
			 | (OP==`BVC_rel & T==`T1BranchCross & phi2)
			 | (OP==`BVC_rel & T==`T1NoBranch & phi2)
			 | (OP==`EOR_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`EOR_izy & T==`Tone & phi2)
			 | (OP==`EOR_izy & T==`Ttwo & phi1)
			 | (OP==`EOR_izy & T==`Tfive & phi2)
			 | (OP==`EOR_zpx & T==`Tone & phi2)
			 | (OP==`EOR_zpx & T==`Ttwo & phi1)
			 | (OP==`LSR_zpx & T==`Tzero & phi1)
			 | (OP==`LSR_zpx & T==`Tone & phi2)
			 | (OP==`LSR_zpx & T==`Ttwo & phi1)
			 | (OP==`LSR_zpx & T==`Tfive & phi2)
			 | (OP==`CLI & T==`Tone & phi2)
			 | (OP==`CLI & T==`Ttwo & phi1)
			 | (OP==`EOR_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`EOR_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`EOR_aby & T==`Tone & phi2)
			 | (OP==`EOR_aby & T==`Ttwo & phi1)
			 | (OP==`EOR_aby & T==`Tfour & phi2)
			 | (OP==`EOR_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`EOR_abx & T==`Tone & phi2)
			 | (OP==`EOR_abx & T==`Ttwo & phi1)
			 | (OP==`EOR_abx & T==`Tfour & phi2)
			 | (OP==`LSR_abx & T==`Tzero & phi1)
			 | (OP==`LSR_abx & T==`Tone & phi2)
			 | (OP==`LSR_abx & T==`Ttwo & phi1)
			 | (OP==`LSR_abx & T==`Tfour & phi2)
			 | (OP==`LSR_abx & T==`Tfive & phi1)
			 | (OP==`LSR_abx & T==`Tsix & phi2)
			 | (OP==`RTS & T==`Tone & phi2)
			 | (OP==`RTS & T==`Ttwo & phi1)
			 | (OP==`RTS & T==`Tfour & phi2)
			 | (OP==`RTS & T==`Tfive & phi1)
			 | (OP==`ADC_izx & T==`Tone & phi2)
			 | (OP==`ADC_izx & T==`Ttwo & phi1)
			 | (OP==`ADC_zp & T==`Tone & phi2)
			 | (OP==`ADC_zp & T==`Ttwo & phi1)
			 | (OP==`ROR_zp & T==`Tzero & phi1)
			 | (OP==`ROR_zp & T==`Tone & phi2)
			 | (OP==`ROR_zp & T==`Ttwo & phi1)
			 | (OP==`ROR_zp & T==`Tfour & phi2)
			 | (OP==`PLA & T==`Tzero & phi1)
			 | (OP==`PLA & T==`Tone & phi2)
			 | (OP==`PLA & T==`Ttwo & phi1)
			 | (OP==`PLA & T==`Tthree & phi2)
			 | (OP==`ADC_imm & T==`Tone & phi2)
			 | (OP==`ADC_imm & T==`Ttwo & phi1)
			 | (OP==`ROR & T==`Tone & phi2)
			 | (OP==`ROR & T==`Ttwo & phi1)
			 | (OP==`JMP_zp & T==`Tone & phi2)
			 | (OP==`JMP_zp & T==`Ttwo & phi1)
			 | (OP==`ADC_abs & T==`Tone & phi2)
			 | (OP==`ADC_abs & T==`Ttwo & phi1)
			 | (OP==`ROR_abs & T==`Tzero & phi1)
			 | (OP==`ROR_abs & T==`Tone & phi2)
			 | (OP==`ROR_abs & T==`Ttwo & phi1)
			 | (OP==`ROR_abs & T==`Tfive & phi2)
			 | (OP==`BVS_rel & T==`Tzero & phi2)
			 | (OP==`BVS_rel & T==`Ttwo & phi1)
			 | (OP==`BVS_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BVS_rel & T==`T1BranchCross & phi1)
			 | (OP==`BVS_rel & T==`T1BranchCross & phi2)
			 | (OP==`BVS_rel & T==`T1NoBranch & phi2)
			 | (OP==`ADC_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`ADC_izy & T==`Tone & phi2)
			 | (OP==`ADC_izy & T==`Ttwo & phi1)
			 | (OP==`ADC_izy & T==`Tfive & phi2)
			 | (OP==`ADC_zpx & T==`Tone & phi2)
			 | (OP==`ADC_zpx & T==`Ttwo & phi1)
			 | (OP==`ROR_zpx & T==`Tzero & phi1)
			 | (OP==`ROR_zpx & T==`Tone & phi2)
			 | (OP==`ROR_zpx & T==`Ttwo & phi1)
			 | (OP==`ROR_zpx & T==`Tfive & phi2)
			 | (OP==`SEI & T==`Tone & phi2)
			 | (OP==`SEI & T==`Ttwo & phi1)
			 | (OP==`ADC_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`ADC_aby & T==`Tone & phi2)
			 | (OP==`ADC_aby & T==`Ttwo & phi1)
			 | (OP==`ADC_aby & T==`Tfour & phi2)
			 | (OP==`ADC_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`ADC_abx & T==`Tone & phi2)
			 | (OP==`ADC_abx & T==`Ttwo & phi1)
			 | (OP==`ADC_abx & T==`Tfour & phi2)
			 | (OP==`ROR_abx & T==`Tzero & phi1)
			 | (OP==`ROR_abx & T==`Tone & phi2)
			 | (OP==`ROR_abx & T==`Ttwo & phi1)
			 | (OP==`ROR_abx & T==`Tfour & phi2)
			 | (OP==`ROR_abx & T==`Tfive & phi1)
			 | (OP==`ROR_abx & T==`Tsix & phi2)
			 | (OP==`STA_izx & T==`Tone & phi2)
			 | (OP==`STA_izx & T==`Ttwo & phi1)
			 | (OP==`STY_zp & T==`Tone & phi2)
			 | (OP==`STY_zp & T==`Ttwo & phi1)
			 | (OP==`STA_zp & T==`Tone & phi2)
			 | (OP==`STA_zp & T==`Ttwo & phi1)
			 | (OP==`STX_zp & T==`Tone & phi2)
			 | (OP==`STX_zp & T==`Ttwo & phi1)
			 | (OP==`DEY & T==`Tone & phi2)
			 | (OP==`DEY & T==`Ttwo & phi1)
			 | (OP==`TXA & T==`Tone & phi2)
			 | (OP==`TXA & T==`Ttwo & phi1)
			 | (OP==`STY_abs & T==`Tone & phi2)
			 | (OP==`STY_abs & T==`Ttwo & phi1)
			 | (OP==`STA_abs & T==`Tone & phi2)
			 | (OP==`STA_abs & T==`Ttwo & phi1)
			 | (OP==`STX_abs & T==`Tone & phi2)
			 | (OP==`STX_abs & T==`Ttwo & phi1)
			 | (OP==`BCC_rel & T==`Tzero & phi2)
			 | (OP==`BCC_rel & T==`Ttwo & phi1)
			 | (OP==`BCC_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BCC_rel & T==`T1BranchCross & phi1)
			 | (OP==`BCC_rel & T==`T1BranchCross & phi2)
			 | (OP==`BCC_rel & T==`T1NoBranch & phi2)
			 | (OP==`STA_izy & T==`Tzero & phi1)
			 | (OP==`STA_izy & T==`Tone & phi2)
			 | (OP==`STA_izy & T==`Ttwo & phi1)
			 | (OP==`STA_izy & T==`Tfive & phi2)
			 | (OP==`STY_zpx & T==`Tone & phi2)
			 | (OP==`STY_zpx & T==`Ttwo & phi1)
			 | (OP==`STA_zpx & T==`Tone & phi2)
			 | (OP==`STA_zpx & T==`Ttwo & phi1)
			 | (OP==`STX_zpy & T==`Tone & phi2)
			 | (OP==`STX_zpy & T==`Ttwo & phi1)
			 | (OP==`TYA & T==`Tone & phi2)
			 | (OP==`TYA & T==`Ttwo & phi1)
			 | (OP==`STA_aby & T==`Tzero & phi1)
			 | (OP==`STA_aby & T==`Tone & phi2)
			 | (OP==`STA_aby & T==`Ttwo & phi1)
			 | (OP==`STA_aby & T==`Tfour & phi2)
			 | (OP==`TXS & T==`Tone & phi2)
			 | (OP==`TXS & T==`Ttwo & phi1)
			 | (OP==`STA_abx & T==`Tzero & phi1)
			 | (OP==`STA_abx & T==`Tone & phi2)
			 | (OP==`STA_abx & T==`Ttwo & phi1)
			 | (OP==`STA_abx & T==`Tfour & phi2)
			 | (OP==`LDY_imm & T==`Tone & phi2)
			 | (OP==`LDY_imm & T==`Ttwo & phi1)
			 | (OP==`LDA_izx & T==`Tone & phi2)
			 | (OP==`LDA_izx & T==`Ttwo & phi1)
			 | (OP==`LDX_imm & T==`Tone & phi2)
			 | (OP==`LDX_imm & T==`Ttwo & phi1)
			 | (OP==`LDY_zp & T==`Tone & phi2)
			 | (OP==`LDY_zp & T==`Ttwo & phi1)
			 | (OP==`LDA_zp & T==`Tone & phi2)
			 | (OP==`LDA_zp & T==`Ttwo & phi1)
			 | (OP==`LDX_zp & T==`Tone & phi2)
			 | (OP==`LDX_zp & T==`Ttwo & phi1)
			 | (OP==`TAY & T==`Tone & phi2)
			 | (OP==`TAY & T==`Ttwo & phi1)
			 | (OP==`LDA_imm & T==`Tone & phi2)
			 | (OP==`LDA_imm & T==`Ttwo & phi1)
			 | (OP==`TAX & T==`Tone & phi2)
			 | (OP==`TAX & T==`Ttwo & phi1)
			 | (OP==`LDY_abs & T==`Tone & phi2)
			 | (OP==`LDY_abs & T==`Ttwo & phi1)
			 | (OP==`LDA_abs & T==`Tone & phi2)
			 | (OP==`LDA_abs & T==`Ttwo & phi1)
			 | (OP==`LDX_abs & T==`Tone & phi2)
			 | (OP==`LDX_abs & T==`Ttwo & phi1)
			 | (OP==`BCS_rel & T==`Tzero & phi2)
			 | (OP==`BCS_rel & T==`Ttwo & phi1)
			 | (OP==`BCS_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BCS_rel & T==`T1BranchCross & phi1)
			 | (OP==`BCS_rel & T==`T1BranchCross & phi2)
			 | (OP==`BCS_rel & T==`T1NoBranch & phi2)
			 | (OP==`LDA_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`LDA_izy & T==`Tone & phi2)
			 | (OP==`LDA_izy & T==`Ttwo & phi1)
			 | (OP==`LDA_izy & T==`Tfive & phi2)
			 | (OP==`LDY_zpx & T==`Tone & phi2)
			 | (OP==`LDY_zpx & T==`Ttwo & phi1)
			 | (OP==`LDA_zpx & T==`Tone & phi2)
			 | (OP==`LDA_zpx & T==`Ttwo & phi1)
			 | (OP==`LDX_zpy & T==`Tone & phi2)
			 | (OP==`LDX_zpy & T==`Ttwo & phi1)
			 | (OP==`CLV & T==`Tone & phi2)
			 | (OP==`CLV & T==`Ttwo & phi1)
			 | (OP==`LDA_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`LDA_aby & T==`Tone & phi2)
			 | (OP==`LDA_aby & T==`Ttwo & phi1)
			 | (OP==`LDA_aby & T==`Tfour & phi2)
			 | (OP==`TSX & T==`Tone & phi2)
			 | (OP==`TSX & T==`Ttwo & phi1)
			 | (OP==`LDY_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`LDY_abx & T==`Tone & phi2)
			 | (OP==`LDY_abx & T==`Ttwo & phi1)
			 | (OP==`LDY_abx & T==`Tfour & phi2)
			 | (OP==`LDA_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`LDA_abx & T==`Tone & phi2)
			 | (OP==`LDA_abx & T==`Ttwo & phi1)
			 | (OP==`LDA_abx & T==`Tfour & phi2)
			 | (OP==`LDX_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`LDX_aby & T==`Tone & phi2)
			 | (OP==`LDX_aby & T==`Ttwo & phi1)
			 | (OP==`LDX_aby & T==`Tfour & phi2)
			 | (OP==`CPY_imm & T==`Tone & phi2)
			 | (OP==`CPY_imm & T==`Ttwo & phi1)
			 | (OP==`CMP_izx & T==`Tone & phi2)
			 | (OP==`CMP_izx & T==`Ttwo & phi1)
			 | (OP==`CPY_zp & T==`Tone & phi2)
			 | (OP==`CPY_zp & T==`Ttwo & phi1)
			 | (OP==`CMP_zp & T==`Tone & phi2)
			 | (OP==`CMP_zp & T==`Ttwo & phi1)
			 | (OP==`DEC_zp & T==`Tzero & phi1)
			 | (OP==`DEC_zp & T==`Tone & phi2)
			 | (OP==`DEC_zp & T==`Ttwo & phi1)
			 | (OP==`DEC_zp & T==`Tfour & phi2)
			 | (OP==`INY & T==`Tone & phi2)
			 | (OP==`INY & T==`Ttwo & phi1)
			 | (OP==`CMP_imm & T==`Tone & phi2)
			 | (OP==`CMP_imm & T==`Ttwo & phi1)
			 | (OP==`DEX & T==`Tone & phi2)
			 | (OP==`DEX & T==`Ttwo & phi1)
			 | (OP==`CPY_abs & T==`Tone & phi2)
			 | (OP==`CPY_abs & T==`Ttwo & phi1)
			 | (OP==`CMP_abs & T==`Tone & phi2)
			 | (OP==`CMP_abs & T==`Ttwo & phi1)
			 | (OP==`DEC_abs & T==`Tzero & phi1)
			 | (OP==`DEC_abs & T==`Tone & phi2)
			 | (OP==`DEC_abs & T==`Ttwo & phi1)
			 | (OP==`DEC_abs & T==`Tfive & phi2)
			 | (OP==`BNE_rel & T==`Tzero & phi2)
			 | (OP==`BNE_rel & T==`Ttwo & phi1)
			 | (OP==`BNE_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BNE_rel & T==`T1BranchCross & phi1)
			 | (OP==`BNE_rel & T==`T1BranchCross & phi2)
			 | (OP==`BNE_rel & T==`T1NoBranch & phi2)
			 | (OP==`CMP_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`CMP_izy & T==`Tone & phi2)
			 | (OP==`CMP_izy & T==`Ttwo & phi1)
			 | (OP==`CMP_izy & T==`Tfive & phi2)
			 | (OP==`CMP_zpx & T==`Tone & phi2)
			 | (OP==`CMP_zpx & T==`Ttwo & phi1)
			 | (OP==`DEC_zpx & T==`Tzero & phi1)
			 | (OP==`DEC_zpx & T==`Tone & phi2)
			 | (OP==`DEC_zpx & T==`Ttwo & phi1)
			 | (OP==`DEC_zpx & T==`Tfive & phi2)
			 | (OP==`CLD & T==`Tone & phi2)
			 | (OP==`CLD & T==`Ttwo & phi1)
			 | (OP==`CMP_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`CMP_aby & T==`Tone & phi2)
			 | (OP==`CMP_aby & T==`Ttwo & phi1)
			 | (OP==`CMP_aby & T==`Tfour & phi2)
			 | (OP==`CMP_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`CMP_abx & T==`Tone & phi2)
			 | (OP==`CMP_abx & T==`Ttwo & phi1)
			 | (OP==`CMP_abx & T==`Tfour & phi2)
			 | (OP==`DEC_abx & T==`Tzero & phi1)
			 | (OP==`DEC_abx & T==`Tone & phi2)
			 | (OP==`DEC_abx & T==`Ttwo & phi1)
			 | (OP==`DEC_abx & T==`Tfour & phi2)
			 | (OP==`DEC_abx & T==`Tfive & phi1)
			 | (OP==`DEC_abx & T==`Tsix & phi2)
			 | (OP==`CPX_imm & T==`Tone & phi2)
			 | (OP==`CPX_imm & T==`Ttwo & phi1)
			 | (OP==`SBC_izx & T==`Tone & phi2)
			 | (OP==`SBC_izx & T==`Ttwo & phi1)
			 | (OP==`CPX_zp & T==`Tone & phi2)
			 | (OP==`CPX_zp & T==`Ttwo & phi1)
			 | (OP==`SBC_zp & T==`Tone & phi2)
			 | (OP==`SBC_zp & T==`Ttwo & phi1)
			 | (OP==`INC_zp & T==`Tzero & phi1)
			 | (OP==`INC_zp & T==`Tone & phi2)
			 | (OP==`INC_zp & T==`Ttwo & phi1)
			 | (OP==`INC_zp & T==`Tfour & phi2)
			 | (OP==`INX & T==`Tone & phi2)
			 | (OP==`INX & T==`Ttwo & phi1)
			 | (OP==`SBC_imm & T==`Tone & phi2)
			 | (OP==`SBC_imm & T==`Ttwo & phi1)
			 | (OP==`NOP & T==`Tone & phi2)
			 | (OP==`NOP & T==`Ttwo & phi1)
			 | (OP==`CPX_abs & T==`Tone & phi2)
			 | (OP==`CPX_abs & T==`Ttwo & phi1)
			 | (OP==`SBC_abs & T==`Tone & phi2)
			 | (OP==`SBC_abs & T==`Ttwo & phi1)
			 | (OP==`INC_abs & T==`Tzero & phi1)
			 | (OP==`INC_abs & T==`Tone & phi2)
			 | (OP==`INC_abs & T==`Ttwo & phi1)
			 | (OP==`INC_abs & T==`Tfive & phi2)
			 | (OP==`BEQ_rel & T==`Tzero & phi2)
			 | (OP==`BEQ_rel & T==`Ttwo & phi1)
			 | (OP==`BEQ_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BEQ_rel & T==`T1BranchCross & phi1)
			 | (OP==`BEQ_rel & T==`T1BranchCross & phi2)
			 | (OP==`BEQ_rel & T==`T1NoBranch & phi2)
			 | (OP==`SBC_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`SBC_izy & T==`Tone & phi2)
			 | (OP==`SBC_izy & T==`Ttwo & phi1)
			 | (OP==`SBC_izy & T==`Tfive & phi2)
			 | (OP==`SBC_zpx & T==`Tone & phi2)
			 | (OP==`SBC_zpx & T==`Ttwo & phi1)
			 | (OP==`INC_zpx & T==`Tzero & phi1)
			 | (OP==`INC_zpx & T==`Tone & phi2)
			 | (OP==`INC_zpx & T==`Ttwo & phi1)
			 | (OP==`INC_zpx & T==`Tfive & phi2)
			 | (OP==`SED & T==`Tone & phi2)
			 | (OP==`SED & T==`Ttwo & phi1)
			 | (OP==`SBC_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`SBC_aby & T==`Tone & phi2)
			 | (OP==`SBC_aby & T==`Ttwo & phi1)
			 | (OP==`SBC_aby & T==`Tfour & phi2)
			 | (OP==`SBC_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`SBC_abx & T==`Tone & phi2)
			 | (OP==`SBC_abx & T==`Ttwo & phi1)
			 | (OP==`SBC_abx & T==`Tfour & phi2)
			 | (OP==`INC_abx & T==`Tzero & phi1)
			 | (OP==`INC_abx & T==`Tone & phi2)
			 | (OP==`INC_abx & T==`Ttwo & phi1)
			 | (OP==`INC_abx & T==`Tfour & phi2)
			 | (OP==`INC_abx & T==`Tfive & phi1)
			 | (OP==`INC_abx & T==`Tsix & phi2)
			;

assign control[`ADD_SB7] = (OP==`BRK & T==`Tone & phi2)
			 | (OP==`BRK & T==`Ttwo & phi1)
			 | (OP==`BRK & T==`Tfive & phi2)
			 | (OP==`BRK & T==`Tsix & phi1)
			 | (OP==`ORA_izx & T==`Tone & phi2)
			 | (OP==`ORA_izx & T==`Ttwo & phi1)
			 | (OP==`ORA_zp & T==`Tone & phi2)
			 | (OP==`ORA_zp & T==`Ttwo & phi1)
			 | (OP==`ASL_zp & T==`Tzero & phi1)
			 | (OP==`ASL_zp & T==`Tone & phi2)
			 | (OP==`ASL_zp & T==`Ttwo & phi1)
			 | (OP==`ASL_zp & T==`Tfour & phi2)
			 | (OP==`PHP & T==`Tzero & phi2)
			 | (OP==`PHP & T==`Tone & phi1)
			 | (OP==`PHP & T==`Tone & phi2)
			 | (OP==`PHP & T==`Ttwo & phi1)
			 | (OP==`ORA_imm & T==`Tone & phi2)
			 | (OP==`ORA_imm & T==`Ttwo & phi1)
			 | (OP==`ASL & T==`Tone & phi2)
			 | (OP==`ASL & T==`Ttwo & phi1)
			 | (OP==`ORA_abs & T==`Tone & phi2)
			 | (OP==`ORA_abs & T==`Ttwo & phi1)
			 | (OP==`ASL_abs & T==`Tzero & phi1)
			 | (OP==`ASL_abs & T==`Tone & phi2)
			 | (OP==`ASL_abs & T==`Ttwo & phi1)
			 | (OP==`ASL_abs & T==`Tfive & phi2)
			 | (OP==`BPL_rel & T==`Tzero & phi2)
			 | (OP==`BPL_rel & T==`Ttwo & phi1)
			 | (OP==`BPL_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BPL_rel & T==`T1BranchCross & phi1)
			 | (OP==`BPL_rel & T==`T1BranchCross & phi2)
			 | (OP==`BPL_rel & T==`T1NoBranch & phi2)
			 | (OP==`ORA_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`ORA_izy & T==`Tone & phi2)
			 | (OP==`ORA_izy & T==`Ttwo & phi1)
			 | (OP==`ORA_izy & T==`Tfive & phi2)
			 | (OP==`ORA_zpx & T==`Tone & phi2)
			 | (OP==`ORA_zpx & T==`Ttwo & phi1)
			 | (OP==`ASL_zpx & T==`Tzero & phi1)
			 | (OP==`ASL_zpx & T==`Tone & phi2)
			 | (OP==`ASL_zpx & T==`Ttwo & phi1)
			 | (OP==`ASL_zpx & T==`Tfive & phi2)
			 | (OP==`CLC & T==`Tone & phi2)
			 | (OP==`CLC & T==`Ttwo & phi1)
			 | (OP==`ORA_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`ORA_aby & T==`Tone & phi2)
			 | (OP==`ORA_aby & T==`Ttwo & phi1)
			 | (OP==`ORA_aby & T==`Tfour & phi2)
			 | (OP==`ORA_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`ORA_abx & T==`Tone & phi2)
			 | (OP==`ORA_abx & T==`Ttwo & phi1)
			 | (OP==`ORA_abx & T==`Tfour & phi2)
			 | (OP==`ASL_abx & T==`Tzero & phi1)
			 | (OP==`ASL_abx & T==`Tone & phi2)
			 | (OP==`ASL_abx & T==`Ttwo & phi1)
			 | (OP==`ASL_abx & T==`Tfour & phi2)
			 | (OP==`ASL_abx & T==`Tfive & phi1)
			 | (OP==`ASL_abx & T==`Tsix & phi2)
			 | (OP==`JSR_abs & T==`Tzero & phi1)
			 | (OP==`JSR_abs & T==`Tzero & phi2)
			 | (OP==`JSR_abs & T==`Tone & phi1)
			 | (OP==`JSR_abs & T==`Tone & phi2)
			 | (OP==`JSR_abs & T==`Ttwo & phi1)
			 | (OP==`JSR_abs & T==`Tfive & phi2)
			 | (OP==`AND_izx & T==`Tone & phi2)
			 | (OP==`AND_izx & T==`Ttwo & phi1)
			 | (OP==`BIT_zp & T==`Tone & phi2)
			 | (OP==`BIT_zp & T==`Ttwo & phi1)
			 | (OP==`AND_zp & T==`Tone & phi2)
			 | (OP==`AND_zp & T==`Ttwo & phi1)
			 | (OP==`ROL_zp & T==`Tzero & phi1)
			 | (OP==`ROL_zp & T==`Tone & phi2)
			 | (OP==`ROL_zp & T==`Ttwo & phi1)
			 | (OP==`ROL_zp & T==`Tfour & phi2)
			 | (OP==`PLP & T==`Tzero & phi1)
			 | (OP==`PLP & T==`Tone & phi2)
			 | (OP==`PLP & T==`Ttwo & phi1)
			 | (OP==`PLP & T==`Tthree & phi2)
			 | (OP==`AND_imm & T==`Tone & phi2)
			 | (OP==`AND_imm & T==`Ttwo & phi1)
			 | (OP==`ROL & T==`Tone & phi2)
			 | (OP==`ROL & T==`Ttwo & phi1)
			 | (OP==`BIT_abs & T==`Tone & phi2)
			 | (OP==`BIT_abs & T==`Ttwo & phi1)
			 | (OP==`AND_abs & T==`Tone & phi2)
			 | (OP==`AND_abs & T==`Ttwo & phi1)
			 | (OP==`ROL_abs & T==`Tzero & phi1)
			 | (OP==`ROL_abs & T==`Tone & phi2)
			 | (OP==`ROL_abs & T==`Ttwo & phi1)
			 | (OP==`ROL_abs & T==`Tfive & phi2)
			 | (OP==`BMI_rel & T==`Tzero & phi2)
			 | (OP==`BMI_rel & T==`Ttwo & phi1)
			 | (OP==`BMI_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BMI_rel & T==`T1BranchCross & phi1)
			 | (OP==`BMI_rel & T==`T1BranchCross & phi2)
			 | (OP==`BMI_rel & T==`T1NoBranch & phi2)
			 | (OP==`AND_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`AND_izy & T==`Tone & phi2)
			 | (OP==`AND_izy & T==`Ttwo & phi1)
			 | (OP==`AND_izy & T==`Tfive & phi2)
			 | (OP==`AND_zpx & T==`Tone & phi2)
			 | (OP==`AND_zpx & T==`Ttwo & phi1)
			 | (OP==`ROL_zpx & T==`Tzero & phi1)
			 | (OP==`ROL_zpx & T==`Tone & phi2)
			 | (OP==`ROL_zpx & T==`Ttwo & phi1)
			 | (OP==`ROL_zpx & T==`Tfive & phi2)
			 | (OP==`SEC & T==`Tone & phi2)
			 | (OP==`SEC & T==`Ttwo & phi1)
			 | (OP==`AND_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`AND_aby & T==`Tone & phi2)
			 | (OP==`AND_aby & T==`Ttwo & phi1)
			 | (OP==`AND_aby & T==`Tfour & phi2)
			 | (OP==`AND_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`AND_abx & T==`Tone & phi2)
			 | (OP==`AND_abx & T==`Ttwo & phi1)
			 | (OP==`AND_abx & T==`Tfour & phi2)
			 | (OP==`ROL_abx & T==`Tzero & phi1)
			 | (OP==`ROL_abx & T==`Tone & phi2)
			 | (OP==`ROL_abx & T==`Ttwo & phi1)
			 | (OP==`ROL_abx & T==`Tfour & phi2)
			 | (OP==`ROL_abx & T==`Tfive & phi1)
			 | (OP==`ROL_abx & T==`Tsix & phi2)
			 | (OP==`RTI & T==`Tzero & phi1)
			 | (OP==`RTI & T==`Tone & phi2)
			 | (OP==`RTI & T==`Ttwo & phi1)
			 | (OP==`RTI & T==`Tfive & phi2)
			 | (OP==`EOR_izx & T==`Tone & phi2)
			 | (OP==`EOR_izx & T==`Ttwo & phi1)
			 | (OP==`EOR_zp & T==`Tone & phi2)
			 | (OP==`EOR_zp & T==`Ttwo & phi1)
			 | (OP==`LSR_zp & T==`Tzero & phi1)
			 | (OP==`LSR_zp & T==`Tone & phi2)
			 | (OP==`LSR_zp & T==`Ttwo & phi1)
			 | (OP==`LSR_zp & T==`Tfour & phi2)
			 | (OP==`PHA & T==`Tzero & phi2)
			 | (OP==`PHA & T==`Tone & phi1)
			 | (OP==`PHA & T==`Tone & phi2)
			 | (OP==`PHA & T==`Ttwo & phi1)
			 | (OP==`EOR_imm & T==`Tone & phi2)
			 | (OP==`EOR_imm & T==`Ttwo & phi1)
			 | (OP==`LSR & T==`Tone & phi2)
			 | (OP==`LSR & T==`Ttwo & phi1)
			 | (OP==`JMP_abs & T==`Tone & phi2)
			 | (OP==`JMP_abs & T==`Ttwo & phi1)
			 | (OP==`EOR_abs & T==`Tone & phi2)
			 | (OP==`EOR_abs & T==`Ttwo & phi1)
			 | (OP==`LSR_abs & T==`Tzero & phi1)
			 | (OP==`LSR_abs & T==`Tone & phi2)
			 | (OP==`LSR_abs & T==`Ttwo & phi1)
			 | (OP==`LSR_abs & T==`Tfive & phi2)
			 | (OP==`BVC_rel & T==`Tzero & phi2)
			 | (OP==`BVC_rel & T==`Ttwo & phi1)
			 | (OP==`BVC_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BVC_rel & T==`T1BranchCross & phi1)
			 | (OP==`BVC_rel & T==`T1BranchCross & phi2)
			 | (OP==`BVC_rel & T==`T1NoBranch & phi2)
			 | (OP==`EOR_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`EOR_izy & T==`Tone & phi2)
			 | (OP==`EOR_izy & T==`Ttwo & phi1)
			 | (OP==`EOR_izy & T==`Tfive & phi2)
			 | (OP==`EOR_zpx & T==`Tone & phi2)
			 | (OP==`EOR_zpx & T==`Ttwo & phi1)
			 | (OP==`LSR_zpx & T==`Tzero & phi1)
			 | (OP==`LSR_zpx & T==`Tone & phi2)
			 | (OP==`LSR_zpx & T==`Ttwo & phi1)
			 | (OP==`LSR_zpx & T==`Tfive & phi2)
			 | (OP==`CLI & T==`Tone & phi2)
			 | (OP==`CLI & T==`Ttwo & phi1)
			 | (OP==`EOR_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`EOR_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`EOR_aby & T==`Tone & phi2)
			 | (OP==`EOR_aby & T==`Ttwo & phi1)
			 | (OP==`EOR_aby & T==`Tfour & phi2)
			 | (OP==`EOR_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`EOR_abx & T==`Tone & phi2)
			 | (OP==`EOR_abx & T==`Ttwo & phi1)
			 | (OP==`EOR_abx & T==`Tfour & phi2)
			 | (OP==`LSR_abx & T==`Tzero & phi1)
			 | (OP==`LSR_abx & T==`Tone & phi2)
			 | (OP==`LSR_abx & T==`Ttwo & phi1)
			 | (OP==`LSR_abx & T==`Tfour & phi2)
			 | (OP==`LSR_abx & T==`Tfive & phi1)
			 | (OP==`LSR_abx & T==`Tsix & phi2)
			 | (OP==`RTS & T==`Tone & phi2)
			 | (OP==`RTS & T==`Ttwo & phi1)
			 | (OP==`RTS & T==`Tfour & phi2)
			 | (OP==`RTS & T==`Tfive & phi1)
			 | (OP==`ADC_izx & T==`Tone & phi2)
			 | (OP==`ADC_izx & T==`Ttwo & phi1)
			 | (OP==`ADC_zp & T==`Tone & phi2)
			 | (OP==`ADC_zp & T==`Ttwo & phi1)
			 | (OP==`ROR_zp & T==`Tzero & phi1)
			 | (OP==`ROR_zp & T==`Tone & phi2)
			 | (OP==`ROR_zp & T==`Ttwo & phi1)
			 | (OP==`ROR_zp & T==`Tfour & phi2)
			 | (OP==`PLA & T==`Tzero & phi1)
			 | (OP==`PLA & T==`Tone & phi2)
			 | (OP==`PLA & T==`Ttwo & phi1)
			 | (OP==`PLA & T==`Tthree & phi2)
			 | (OP==`ADC_imm & T==`Tone & phi2)
			 | (OP==`ADC_imm & T==`Ttwo & phi1)
			 | (OP==`ROR & T==`Tone & phi2)
			 | (OP==`ROR & T==`Ttwo & phi1)
			 | (OP==`JMP_zp & T==`Tone & phi2)
			 | (OP==`JMP_zp & T==`Ttwo & phi1)
			 | (OP==`ADC_abs & T==`Tone & phi2)
			 | (OP==`ADC_abs & T==`Ttwo & phi1)
			 | (OP==`ROR_abs & T==`Tzero & phi1)
			 | (OP==`ROR_abs & T==`Tone & phi2)
			 | (OP==`ROR_abs & T==`Ttwo & phi1)
			 | (OP==`ROR_abs & T==`Tfive & phi2)
			 | (OP==`BVS_rel & T==`Tzero & phi2)
			 | (OP==`BVS_rel & T==`Ttwo & phi1)
			 | (OP==`BVS_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BVS_rel & T==`T1BranchCross & phi1)
			 | (OP==`BVS_rel & T==`T1BranchCross & phi2)
			 | (OP==`BVS_rel & T==`T1NoBranch & phi2)
			 | (OP==`ADC_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`ADC_izy & T==`Tone & phi2)
			 | (OP==`ADC_izy & T==`Ttwo & phi1)
			 | (OP==`ADC_izy & T==`Tfive & phi2)
			 | (OP==`ADC_zpx & T==`Tone & phi2)
			 | (OP==`ADC_zpx & T==`Ttwo & phi1)
			 | (OP==`ROR_zpx & T==`Tzero & phi1)
			 | (OP==`ROR_zpx & T==`Tone & phi2)
			 | (OP==`ROR_zpx & T==`Ttwo & phi1)
			 | (OP==`ROR_zpx & T==`Tfive & phi2)
			 | (OP==`SEI & T==`Tone & phi2)
			 | (OP==`SEI & T==`Ttwo & phi1)
			 | (OP==`ADC_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`ADC_aby & T==`Tone & phi2)
			 | (OP==`ADC_aby & T==`Ttwo & phi1)
			 | (OP==`ADC_aby & T==`Tfour & phi2)
			 | (OP==`ADC_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`ADC_abx & T==`Tone & phi2)
			 | (OP==`ADC_abx & T==`Ttwo & phi1)
			 | (OP==`ADC_abx & T==`Tfour & phi2)
			 | (OP==`ROR_abx & T==`Tzero & phi1)
			 | (OP==`ROR_abx & T==`Tone & phi2)
			 | (OP==`ROR_abx & T==`Ttwo & phi1)
			 | (OP==`ROR_abx & T==`Tfour & phi2)
			 | (OP==`ROR_abx & T==`Tfive & phi1)
			 | (OP==`ROR_abx & T==`Tsix & phi2)
			 | (OP==`STA_izx & T==`Tone & phi2)
			 | (OP==`STA_izx & T==`Ttwo & phi1)
			 | (OP==`STY_zp & T==`Tone & phi2)
			 | (OP==`STY_zp & T==`Ttwo & phi1)
			 | (OP==`STA_zp & T==`Tone & phi2)
			 | (OP==`STA_zp & T==`Ttwo & phi1)
			 | (OP==`STX_zp & T==`Tone & phi2)
			 | (OP==`STX_zp & T==`Ttwo & phi1)
			 | (OP==`DEY & T==`Tone & phi2)
			 | (OP==`DEY & T==`Ttwo & phi1)
			 | (OP==`TXA & T==`Tone & phi2)
			 | (OP==`TXA & T==`Ttwo & phi1)
			 | (OP==`STY_abs & T==`Tone & phi2)
			 | (OP==`STY_abs & T==`Ttwo & phi1)
			 | (OP==`STA_abs & T==`Tone & phi2)
			 | (OP==`STA_abs & T==`Ttwo & phi1)
			 | (OP==`STX_abs & T==`Tone & phi2)
			 | (OP==`STX_abs & T==`Ttwo & phi1)
			 | (OP==`BCC_rel & T==`Tzero & phi2)
			 | (OP==`BCC_rel & T==`Ttwo & phi1)
			 | (OP==`BCC_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BCC_rel & T==`T1BranchCross & phi1)
			 | (OP==`BCC_rel & T==`T1BranchCross & phi2)
			 | (OP==`BCC_rel & T==`T1NoBranch & phi2)
			 | (OP==`STA_izy & T==`Tzero & phi1)
			 | (OP==`STA_izy & T==`Tone & phi2)
			 | (OP==`STA_izy & T==`Ttwo & phi1)
			 | (OP==`STA_izy & T==`Tfive & phi2)
			 | (OP==`STY_zpx & T==`Tone & phi2)
			 | (OP==`STY_zpx & T==`Ttwo & phi1)
			 | (OP==`STA_zpx & T==`Tone & phi2)
			 | (OP==`STA_zpx & T==`Ttwo & phi1)
			 | (OP==`STX_zpy & T==`Tone & phi2)
			 | (OP==`STX_zpy & T==`Ttwo & phi1)
			 | (OP==`TYA & T==`Tone & phi2)
			 | (OP==`TYA & T==`Ttwo & phi1)
			 | (OP==`STA_aby & T==`Tzero & phi1)
			 | (OP==`STA_aby & T==`Tone & phi2)
			 | (OP==`STA_aby & T==`Ttwo & phi1)
			 | (OP==`STA_aby & T==`Tfour & phi2)
			 | (OP==`TXS & T==`Tone & phi2)
			 | (OP==`TXS & T==`Ttwo & phi1)
			 | (OP==`STA_abx & T==`Tzero & phi1)
			 | (OP==`STA_abx & T==`Tone & phi2)
			 | (OP==`STA_abx & T==`Ttwo & phi1)
			 | (OP==`STA_abx & T==`Tfour & phi2)
			 | (OP==`LDY_imm & T==`Tone & phi2)
			 | (OP==`LDY_imm & T==`Ttwo & phi1)
			 | (OP==`LDA_izx & T==`Tone & phi2)
			 | (OP==`LDA_izx & T==`Ttwo & phi1)
			 | (OP==`LDX_imm & T==`Tone & phi2)
			 | (OP==`LDX_imm & T==`Ttwo & phi1)
			 | (OP==`LDY_zp & T==`Tone & phi2)
			 | (OP==`LDY_zp & T==`Ttwo & phi1)
			 | (OP==`LDA_zp & T==`Tone & phi2)
			 | (OP==`LDA_zp & T==`Ttwo & phi1)
			 | (OP==`LDX_zp & T==`Tone & phi2)
			 | (OP==`LDX_zp & T==`Ttwo & phi1)
			 | (OP==`TAY & T==`Tone & phi2)
			 | (OP==`TAY & T==`Ttwo & phi1)
			 | (OP==`LDA_imm & T==`Tone & phi2)
			 | (OP==`LDA_imm & T==`Ttwo & phi1)
			 | (OP==`TAX & T==`Tone & phi2)
			 | (OP==`TAX & T==`Ttwo & phi1)
			 | (OP==`LDY_abs & T==`Tone & phi2)
			 | (OP==`LDY_abs & T==`Ttwo & phi1)
			 | (OP==`LDA_abs & T==`Tone & phi2)
			 | (OP==`LDA_abs & T==`Ttwo & phi1)
			 | (OP==`LDX_abs & T==`Tone & phi2)
			 | (OP==`LDX_abs & T==`Ttwo & phi1)
			 | (OP==`BCS_rel & T==`Tzero & phi2)
			 | (OP==`BCS_rel & T==`Ttwo & phi1)
			 | (OP==`BCS_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BCS_rel & T==`T1BranchCross & phi1)
			 | (OP==`BCS_rel & T==`T1BranchCross & phi2)
			 | (OP==`BCS_rel & T==`T1NoBranch & phi2)
			 | (OP==`LDA_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`LDA_izy & T==`Tone & phi2)
			 | (OP==`LDA_izy & T==`Ttwo & phi1)
			 | (OP==`LDA_izy & T==`Tfive & phi2)
			 | (OP==`LDY_zpx & T==`Tone & phi2)
			 | (OP==`LDY_zpx & T==`Ttwo & phi1)
			 | (OP==`LDA_zpx & T==`Tone & phi2)
			 | (OP==`LDA_zpx & T==`Ttwo & phi1)
			 | (OP==`LDX_zpy & T==`Tone & phi2)
			 | (OP==`LDX_zpy & T==`Ttwo & phi1)
			 | (OP==`CLV & T==`Tone & phi2)
			 | (OP==`CLV & T==`Ttwo & phi1)
			 | (OP==`LDA_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`LDA_aby & T==`Tone & phi2)
			 | (OP==`LDA_aby & T==`Ttwo & phi1)
			 | (OP==`LDA_aby & T==`Tfour & phi2)
			 | (OP==`TSX & T==`Tone & phi2)
			 | (OP==`TSX & T==`Ttwo & phi1)
			 | (OP==`LDY_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`LDY_abx & T==`Tone & phi2)
			 | (OP==`LDY_abx & T==`Ttwo & phi1)
			 | (OP==`LDY_abx & T==`Tfour & phi2)
			 | (OP==`LDA_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`LDA_abx & T==`Tone & phi2)
			 | (OP==`LDA_abx & T==`Ttwo & phi1)
			 | (OP==`LDA_abx & T==`Tfour & phi2)
			 | (OP==`LDX_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`LDX_aby & T==`Tone & phi2)
			 | (OP==`LDX_aby & T==`Ttwo & phi1)
			 | (OP==`LDX_aby & T==`Tfour & phi2)
			 | (OP==`CPY_imm & T==`Tone & phi2)
			 | (OP==`CPY_imm & T==`Ttwo & phi1)
			 | (OP==`CMP_izx & T==`Tone & phi2)
			 | (OP==`CMP_izx & T==`Ttwo & phi1)
			 | (OP==`CPY_zp & T==`Tone & phi2)
			 | (OP==`CPY_zp & T==`Ttwo & phi1)
			 | (OP==`CMP_zp & T==`Tone & phi2)
			 | (OP==`CMP_zp & T==`Ttwo & phi1)
			 | (OP==`DEC_zp & T==`Tzero & phi1)
			 | (OP==`DEC_zp & T==`Tone & phi2)
			 | (OP==`DEC_zp & T==`Ttwo & phi1)
			 | (OP==`DEC_zp & T==`Tfour & phi2)
			 | (OP==`INY & T==`Tone & phi2)
			 | (OP==`INY & T==`Ttwo & phi1)
			 | (OP==`CMP_imm & T==`Tone & phi2)
			 | (OP==`CMP_imm & T==`Ttwo & phi1)
			 | (OP==`DEX & T==`Tone & phi2)
			 | (OP==`DEX & T==`Ttwo & phi1)
			 | (OP==`CPY_abs & T==`Tone & phi2)
			 | (OP==`CPY_abs & T==`Ttwo & phi1)
			 | (OP==`CMP_abs & T==`Tone & phi2)
			 | (OP==`CMP_abs & T==`Ttwo & phi1)
			 | (OP==`DEC_abs & T==`Tzero & phi1)
			 | (OP==`DEC_abs & T==`Tone & phi2)
			 | (OP==`DEC_abs & T==`Ttwo & phi1)
			 | (OP==`DEC_abs & T==`Tfive & phi2)
			 | (OP==`BNE_rel & T==`Tzero & phi2)
			 | (OP==`BNE_rel & T==`Ttwo & phi1)
			 | (OP==`BNE_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BNE_rel & T==`T1BranchCross & phi1)
			 | (OP==`BNE_rel & T==`T1BranchCross & phi2)
			 | (OP==`BNE_rel & T==`T1NoBranch & phi2)
			 | (OP==`CMP_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`CMP_izy & T==`Tone & phi2)
			 | (OP==`CMP_izy & T==`Ttwo & phi1)
			 | (OP==`CMP_izy & T==`Tfive & phi2)
			 | (OP==`CMP_zpx & T==`Tone & phi2)
			 | (OP==`CMP_zpx & T==`Ttwo & phi1)
			 | (OP==`DEC_zpx & T==`Tzero & phi1)
			 | (OP==`DEC_zpx & T==`Tone & phi2)
			 | (OP==`DEC_zpx & T==`Ttwo & phi1)
			 | (OP==`DEC_zpx & T==`Tfive & phi2)
			 | (OP==`CLD & T==`Tone & phi2)
			 | (OP==`CLD & T==`Ttwo & phi1)
			 | (OP==`CMP_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`CMP_aby & T==`Tone & phi2)
			 | (OP==`CMP_aby & T==`Ttwo & phi1)
			 | (OP==`CMP_aby & T==`Tfour & phi2)
			 | (OP==`CMP_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`CMP_abx & T==`Tone & phi2)
			 | (OP==`CMP_abx & T==`Ttwo & phi1)
			 | (OP==`CMP_abx & T==`Tfour & phi2)
			 | (OP==`DEC_abx & T==`Tzero & phi1)
			 | (OP==`DEC_abx & T==`Tone & phi2)
			 | (OP==`DEC_abx & T==`Ttwo & phi1)
			 | (OP==`DEC_abx & T==`Tfour & phi2)
			 | (OP==`DEC_abx & T==`Tfive & phi1)
			 | (OP==`DEC_abx & T==`Tsix & phi2)
			 | (OP==`CPX_imm & T==`Tone & phi2)
			 | (OP==`CPX_imm & T==`Ttwo & phi1)
			 | (OP==`SBC_izx & T==`Tone & phi2)
			 | (OP==`SBC_izx & T==`Ttwo & phi1)
			 | (OP==`CPX_zp & T==`Tone & phi2)
			 | (OP==`CPX_zp & T==`Ttwo & phi1)
			 | (OP==`SBC_zp & T==`Tone & phi2)
			 | (OP==`SBC_zp & T==`Ttwo & phi1)
			 | (OP==`INC_zp & T==`Tzero & phi1)
			 | (OP==`INC_zp & T==`Tone & phi2)
			 | (OP==`INC_zp & T==`Ttwo & phi1)
			 | (OP==`INC_zp & T==`Tfour & phi2)
			 | (OP==`INX & T==`Tone & phi2)
			 | (OP==`INX & T==`Ttwo & phi1)
			 | (OP==`SBC_imm & T==`Tone & phi2)
			 | (OP==`SBC_imm & T==`Ttwo & phi1)
			 | (OP==`NOP & T==`Tone & phi2)
			 | (OP==`NOP & T==`Ttwo & phi1)
			 | (OP==`CPX_abs & T==`Tone & phi2)
			 | (OP==`CPX_abs & T==`Ttwo & phi1)
			 | (OP==`SBC_abs & T==`Tone & phi2)
			 | (OP==`SBC_abs & T==`Ttwo & phi1)
			 | (OP==`INC_abs & T==`Tzero & phi1)
			 | (OP==`INC_abs & T==`Tone & phi2)
			 | (OP==`INC_abs & T==`Ttwo & phi1)
			 | (OP==`INC_abs & T==`Tfive & phi2)
			 | (OP==`BEQ_rel & T==`Tzero & phi2)
			 | (OP==`BEQ_rel & T==`Ttwo & phi1)
			 | (OP==`BEQ_rel & T==`T1BranchNoCross & phi2)
			 | (OP==`BEQ_rel & T==`T1BranchCross & phi1)
			 | (OP==`BEQ_rel & T==`T1BranchCross & phi2)
			 | (OP==`BEQ_rel & T==`T1NoBranch & phi2)
			 | (OP==`SBC_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`SBC_izy & T==`Tone & phi2)
			 | (OP==`SBC_izy & T==`Ttwo & phi1)
			 | (OP==`SBC_izy & T==`Tfive & phi2)
			 | (OP==`SBC_zpx & T==`Tone & phi2)
			 | (OP==`SBC_zpx & T==`Ttwo & phi1)
			 | (OP==`INC_zpx & T==`Tzero & phi1)
			 | (OP==`INC_zpx & T==`Tone & phi2)
			 | (OP==`INC_zpx & T==`Ttwo & phi1)
			 | (OP==`INC_zpx & T==`Tfive & phi2)
			 | (OP==`SED & T==`Tone & phi2)
			 | (OP==`SED & T==`Ttwo & phi1)
			 | (OP==`SBC_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`SBC_aby & T==`Tone & phi2)
			 | (OP==`SBC_aby & T==`Ttwo & phi1)
			 | (OP==`SBC_aby & T==`Tfour & phi2)
			 | (OP==`SBC_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`SBC_abx & T==`Tone & phi2)
			 | (OP==`SBC_abx & T==`Ttwo & phi1)
			 | (OP==`SBC_abx & T==`Tfour & phi2)
			 | (OP==`INC_abx & T==`Tzero & phi1)
			 | (OP==`INC_abx & T==`Tone & phi2)
			 | (OP==`INC_abx & T==`Ttwo & phi1)
			 | (OP==`INC_abx & T==`Tfour & phi2)
			 | (OP==`INC_abx & T==`Tfive & phi1)
			 | (OP==`INC_abx & T==`Tsix & phi2)
			;

assign control[`O_ADD] = (OP==`BRK & T==`Tzero & phi1)
			 | (OP==`BRK & T==`Tsix & phi1)
			 | (OP==`ORA_izx & T==`Tfour & phi1)
			 | (OP==`ORA_izx & T==`Tfive & phi1)
			 | (OP==`PHP & T==`Tone & phi1)
			 | (OP==`ORA_abs & T==`Tthree & phi1)
			 | (OP==`ASL_abs & T==`Tthree & phi1)
			 | (OP==`ORA_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ORA_izy & T==`Tthree & phi1)
			 | (OP==`ORA_izy & T==`Tfive & phi1)
			 | (OP==`ORA_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ORA_aby & T==`Tfour & phi1)
			 | (OP==`ORA_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ORA_abx & T==`Tfour & phi1)
			 | (OP==`ASL_abx & T==`Tfour & phi1)
			 | (OP==`JSR_abs & T==`Tone & phi1)
			 | (OP==`JSR_abs & T==`Tthree & phi1)
			 | (OP==`AND_izx & T==`Tfour & phi1)
			 | (OP==`AND_izx & T==`Tfive & phi1)
			 | (OP==`PLP & T==`Tzero & phi1)
			 | (OP==`PLP & T==`Tone & phi1)
			 | (OP==`PLP & T==`Tthree & phi1)
			 | (OP==`BIT_abs & T==`Tthree & phi1)
			 | (OP==`AND_abs & T==`Tthree & phi1)
			 | (OP==`ROL_abs & T==`Tthree & phi1)
			 | (OP==`AND_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`AND_izy & T==`Tthree & phi1)
			 | (OP==`AND_izy & T==`Tfive & phi1)
			 | (OP==`AND_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`AND_aby & T==`Tfour & phi1)
			 | (OP==`AND_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`AND_abx & T==`Tfour & phi1)
			 | (OP==`ROL_abx & T==`Tfour & phi1)
			 | (OP==`RTI & T==`Tzero & phi1)
			 | (OP==`RTI & T==`Tone & phi1)
			 | (OP==`RTI & T==`Tthree & phi1)
			 | (OP==`RTI & T==`Tfour & phi1)
			 | (OP==`RTI & T==`Tfive & phi1)
			 | (OP==`EOR_izx & T==`Tfour & phi1)
			 | (OP==`EOR_izx & T==`Tfive & phi1)
			 | (OP==`PHA & T==`Tone & phi1)
			 | (OP==`JMP_abs & T==`Tzero & phi1)
			 | (OP==`JMP_abs & T==`Tone & phi1)
			 | (OP==`EOR_abs & T==`Tthree & phi1)
			 | (OP==`LSR_abs & T==`Tthree & phi1)
			 | (OP==`EOR_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`EOR_izy & T==`Tthree & phi1)
			 | (OP==`EOR_izy & T==`Tfive & phi1)
			 | (OP==`EOR_aby & T==`Tfour & phi1)
			 | (OP==`EOR_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`EOR_abx & T==`Tfour & phi1)
			 | (OP==`LSR_abx & T==`Tfour & phi1)
			 | (OP==`RTS & T==`Tzero & phi1)
			 | (OP==`RTS & T==`Tone & phi1)
			 | (OP==`RTS & T==`Tthree & phi1)
			 | (OP==`RTS & T==`Tfour & phi1)
			 | (OP==`RTS & T==`Tfive & phi1)
			 | (OP==`ADC_izx & T==`Tfour & phi1)
			 | (OP==`ADC_izx & T==`Tfive & phi1)
			 | (OP==`PLA & T==`Tzero & phi1)
			 | (OP==`PLA & T==`Tone & phi1)
			 | (OP==`PLA & T==`Tthree & phi1)
			 | (OP==`JMP_zp & T==`Tzero & phi1)
			 | (OP==`JMP_zp & T==`Tone & phi1)
			 | (OP==`JMP_zp & T==`Tthree & phi1)
			 | (OP==`JMP_zp & T==`Tfour & phi1)
			 | (OP==`ADC_abs & T==`Tthree & phi1)
			 | (OP==`ROR_abs & T==`Tthree & phi1)
			 | (OP==`ADC_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ADC_izy & T==`Tthree & phi1)
			 | (OP==`ADC_izy & T==`Tfive & phi1)
			 | (OP==`ADC_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ADC_aby & T==`Tfour & phi1)
			 | (OP==`ADC_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`ADC_abx & T==`Tfour & phi1)
			 | (OP==`ROR_abx & T==`Tfour & phi1)
			 | (OP==`STA_izx & T==`Tfour & phi1)
			 | (OP==`STA_izx & T==`Tfive & phi1)
			 | (OP==`STY_abs & T==`Tthree & phi1)
			 | (OP==`STA_abs & T==`Tthree & phi1)
			 | (OP==`STX_abs & T==`Tthree & phi1)
			 | (OP==`STA_izy & T==`Tthree & phi1)
			 | (OP==`STA_izy & T==`Tfive & phi1)
			 | (OP==`STA_aby & T==`Tfour & phi1)
			 | (OP==`STA_abx & T==`Tfour & phi1)
			 | (OP==`LDA_izx & T==`Tfour & phi1)
			 | (OP==`LDA_izx & T==`Tfive & phi1)
			 | (OP==`LDY_abs & T==`Tthree & phi1)
			 | (OP==`LDA_abs & T==`Tthree & phi1)
			 | (OP==`LDX_abs & T==`Tthree & phi1)
			 | (OP==`LDA_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDA_izy & T==`Tthree & phi1)
			 | (OP==`LDA_izy & T==`Tfive & phi1)
			 | (OP==`LDA_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDA_aby & T==`Tfour & phi1)
			 | (OP==`LDY_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDY_abx & T==`Tfour & phi1)
			 | (OP==`LDA_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDA_abx & T==`Tfour & phi1)
			 | (OP==`LDX_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`LDX_aby & T==`Tfour & phi1)
			 | (OP==`CMP_izx & T==`Tfour & phi1)
			 | (OP==`CMP_izx & T==`Tfive & phi1)
			 | (OP==`CPY_abs & T==`Tthree & phi1)
			 | (OP==`CMP_abs & T==`Tthree & phi1)
			 | (OP==`DEC_abs & T==`Tthree & phi1)
			 | (OP==`CMP_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`CMP_izy & T==`Tthree & phi1)
			 | (OP==`CMP_izy & T==`Tfive & phi1)
			 | (OP==`CMP_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`CMP_aby & T==`Tfour & phi1)
			 | (OP==`CMP_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`CMP_abx & T==`Tfour & phi1)
			 | (OP==`DEC_abx & T==`Tfour & phi1)
			 | (OP==`SBC_izx & T==`Tfour & phi1)
			 | (OP==`SBC_izx & T==`Tfive & phi1)
			 | (OP==`INC_zp & T==`Tfour & phi1)
			 | (OP==`CPX_abs & T==`Tthree & phi1)
			 | (OP==`SBC_abs & T==`Tthree & phi1)
			 | (OP==`INC_abs & T==`Tthree & phi1)
			 | (OP==`INC_abs & T==`Tfive & phi1)
			 | (OP==`SBC_izy & T==`TzeroNoCrossPg & phi1)
			 | (OP==`SBC_izy & T==`Tthree & phi1)
			 | (OP==`SBC_izy & T==`Tfive & phi1)
			 | (OP==`INC_zpx & T==`Tfive & phi1)
			 | (OP==`SBC_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`SBC_aby & T==`Tfour & phi1)
			 | (OP==`SBC_abx & T==`TzeroNoCrossPg & phi1)
			 | (OP==`SBC_abx & T==`Tfour & phi1)
			 | (OP==`INC_abx & T==`Tfour & phi1)
			 | (OP==`INC_abx & T==`Tsix & phi1)
			;

assign control[`SB_ADD] = (OP==`BRK & T==`Tone & phi1)
			 | (OP==`BRK & T==`Ttwo & phi1)
			 | (OP==`BRK & T==`Tthree & phi1)
			 | (OP==`BRK & T==`Tfour & phi1)
			 | (OP==`BRK & T==`Tfive & phi1)
			 | (OP==`ORA_izx & T==`Tzero & phi1)
			 | (OP==`ORA_izx & T==`Tone & phi1)
			 | (OP==`ORA_izx & T==`Ttwo & phi1)
			 | (OP==`ORA_izx & T==`Tthree & phi1)
			 | (OP==`ORA_zp & T==`Tzero & phi1)
			 | (OP==`ORA_zp & T==`Tone & phi1)
			 | (OP==`ORA_zp & T==`Ttwo & phi1)
			 | (OP==`ASL_zp & T==`Tzero & phi1)
			 | (OP==`ASL_zp & T==`Tone & phi1)
			 | (OP==`ASL_zp & T==`Ttwo & phi1)
			 | (OP==`ASL_zp & T==`Tthree & phi1)
			 | (OP==`ASL_zp & T==`Tfour & phi1)
			 | (OP==`PHP & T==`Tzero & phi1)
			 | (OP==`PHP & T==`Ttwo & phi1)
			 | (OP==`ORA_imm & T==`Tone & phi1)
			 | (OP==`ORA_imm & T==`Ttwo & phi1)
			 | (OP==`ASL & T==`Tone & phi1)
			 | (OP==`ASL & T==`Ttwo & phi1)
			 | (OP==`ORA_abs & T==`Tzero & phi1)
			 | (OP==`ORA_abs & T==`Tone & phi1)
			 | (OP==`ORA_abs & T==`Ttwo & phi1)
			 | (OP==`ASL_abs & T==`Tzero & phi1)
			 | (OP==`ASL_abs & T==`Tone & phi1)
			 | (OP==`ASL_abs & T==`Ttwo & phi1)
			 | (OP==`ASL_abs & T==`Tfour & phi1)
			 | (OP==`ASL_abs & T==`Tfive & phi1)
			 | (OP==`BPL_rel & T==`Tzero & phi1)
			 | (OP==`BPL_rel & T==`Ttwo & phi1)
			 | (OP==`BPL_rel & T==`Tthree & phi1)
			 | (OP==`BPL_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BPL_rel & T==`T1BranchCross & phi1)
			 | (OP==`BPL_rel & T==`T1NoBranch & phi1)
			 | (OP==`ORA_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`ORA_izy & T==`Tone & phi1)
			 | (OP==`ORA_izy & T==`Ttwo & phi1)
			 | (OP==`ORA_izy & T==`Tfour & phi1)
			 | (OP==`ORA_zpx & T==`Tzero & phi1)
			 | (OP==`ORA_zpx & T==`Tone & phi1)
			 | (OP==`ORA_zpx & T==`Ttwo & phi1)
			 | (OP==`ORA_zpx & T==`Tthree & phi1)
			 | (OP==`ASL_zpx & T==`Tzero & phi1)
			 | (OP==`ASL_zpx & T==`Tone & phi1)
			 | (OP==`ASL_zpx & T==`Ttwo & phi1)
			 | (OP==`ASL_zpx & T==`Tthree & phi1)
			 | (OP==`ASL_zpx & T==`Tfour & phi1)
			 | (OP==`ASL_zpx & T==`Tfive & phi1)
			 | (OP==`CLC & T==`Tone & phi1)
			 | (OP==`CLC & T==`Ttwo & phi1)
			 | (OP==`ORA_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`ORA_aby & T==`Tone & phi1)
			 | (OP==`ORA_aby & T==`Ttwo & phi1)
			 | (OP==`ORA_aby & T==`Tthree & phi1)
			 | (OP==`ORA_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`ORA_abx & T==`Tone & phi1)
			 | (OP==`ORA_abx & T==`Ttwo & phi1)
			 | (OP==`ORA_abx & T==`Tthree & phi1)
			 | (OP==`ASL_abx & T==`Tzero & phi1)
			 | (OP==`ASL_abx & T==`Tone & phi1)
			 | (OP==`ASL_abx & T==`Ttwo & phi1)
			 | (OP==`ASL_abx & T==`Tthree & phi1)
			 | (OP==`ASL_abx & T==`Tfive & phi1)
			 | (OP==`ASL_abx & T==`Tsix & phi1)
			 | (OP==`JSR_abs & T==`Tzero & phi1)
			 | (OP==`JSR_abs & T==`Ttwo & phi1)
			 | (OP==`JSR_abs & T==`Tfour & phi1)
			 | (OP==`JSR_abs & T==`Tfive & phi1)
			 | (OP==`AND_izx & T==`Tzero & phi1)
			 | (OP==`AND_izx & T==`Tone & phi1)
			 | (OP==`AND_izx & T==`Ttwo & phi1)
			 | (OP==`AND_izx & T==`Tthree & phi1)
			 | (OP==`BIT_zp & T==`Tzero & phi1)
			 | (OP==`BIT_zp & T==`Tone & phi1)
			 | (OP==`BIT_zp & T==`Ttwo & phi1)
			 | (OP==`AND_zp & T==`Tzero & phi1)
			 | (OP==`AND_zp & T==`Tone & phi1)
			 | (OP==`AND_zp & T==`Ttwo & phi1)
			 | (OP==`ROL_zp & T==`Tzero & phi1)
			 | (OP==`ROL_zp & T==`Tone & phi1)
			 | (OP==`ROL_zp & T==`Ttwo & phi1)
			 | (OP==`ROL_zp & T==`Tthree & phi1)
			 | (OP==`ROL_zp & T==`Tfour & phi1)
			 | (OP==`PLP & T==`Ttwo & phi1)
			 | (OP==`AND_imm & T==`Tone & phi1)
			 | (OP==`AND_imm & T==`Ttwo & phi1)
			 | (OP==`ROL & T==`Tone & phi1)
			 | (OP==`ROL & T==`Ttwo & phi1)
			 | (OP==`BIT_abs & T==`Tzero & phi1)
			 | (OP==`BIT_abs & T==`Tone & phi1)
			 | (OP==`BIT_abs & T==`Ttwo & phi1)
			 | (OP==`AND_abs & T==`Tzero & phi1)
			 | (OP==`AND_abs & T==`Tone & phi1)
			 | (OP==`AND_abs & T==`Ttwo & phi1)
			 | (OP==`ROL_abs & T==`Tzero & phi1)
			 | (OP==`ROL_abs & T==`Tone & phi1)
			 | (OP==`ROL_abs & T==`Ttwo & phi1)
			 | (OP==`ROL_abs & T==`Tfour & phi1)
			 | (OP==`ROL_abs & T==`Tfive & phi1)
			 | (OP==`BMI_rel & T==`Tzero & phi1)
			 | (OP==`BMI_rel & T==`Ttwo & phi1)
			 | (OP==`BMI_rel & T==`Tthree & phi1)
			 | (OP==`BMI_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BMI_rel & T==`T1BranchCross & phi1)
			 | (OP==`BMI_rel & T==`T1NoBranch & phi1)
			 | (OP==`AND_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`AND_izy & T==`Tone & phi1)
			 | (OP==`AND_izy & T==`Ttwo & phi1)
			 | (OP==`AND_izy & T==`Tfour & phi1)
			 | (OP==`AND_zpx & T==`Tzero & phi1)
			 | (OP==`AND_zpx & T==`Tone & phi1)
			 | (OP==`AND_zpx & T==`Ttwo & phi1)
			 | (OP==`AND_zpx & T==`Tthree & phi1)
			 | (OP==`ROL_zpx & T==`Tzero & phi1)
			 | (OP==`ROL_zpx & T==`Tone & phi1)
			 | (OP==`ROL_zpx & T==`Ttwo & phi1)
			 | (OP==`ROL_zpx & T==`Tthree & phi1)
			 | (OP==`ROL_zpx & T==`Tfour & phi1)
			 | (OP==`ROL_zpx & T==`Tfive & phi1)
			 | (OP==`SEC & T==`Tone & phi1)
			 | (OP==`SEC & T==`Ttwo & phi1)
			 | (OP==`AND_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`AND_aby & T==`Tone & phi1)
			 | (OP==`AND_aby & T==`Ttwo & phi1)
			 | (OP==`AND_aby & T==`Tthree & phi1)
			 | (OP==`AND_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`AND_abx & T==`Tone & phi1)
			 | (OP==`AND_abx & T==`Ttwo & phi1)
			 | (OP==`AND_abx & T==`Tthree & phi1)
			 | (OP==`ROL_abx & T==`Tzero & phi1)
			 | (OP==`ROL_abx & T==`Tone & phi1)
			 | (OP==`ROL_abx & T==`Ttwo & phi1)
			 | (OP==`ROL_abx & T==`Tthree & phi1)
			 | (OP==`ROL_abx & T==`Tfive & phi1)
			 | (OP==`ROL_abx & T==`Tsix & phi1)
			 | (OP==`RTI & T==`Ttwo & phi1)
			 | (OP==`EOR_izx & T==`Tzero & phi1)
			 | (OP==`EOR_izx & T==`Tone & phi1)
			 | (OP==`EOR_izx & T==`Ttwo & phi1)
			 | (OP==`EOR_izx & T==`Tthree & phi1)
			 | (OP==`EOR_zp & T==`Tzero & phi1)
			 | (OP==`EOR_zp & T==`Tone & phi1)
			 | (OP==`EOR_zp & T==`Ttwo & phi1)
			 | (OP==`LSR_zp & T==`Tzero & phi1)
			 | (OP==`LSR_zp & T==`Tone & phi1)
			 | (OP==`LSR_zp & T==`Ttwo & phi1)
			 | (OP==`LSR_zp & T==`Tthree & phi1)
			 | (OP==`LSR_zp & T==`Tfour & phi1)
			 | (OP==`PHA & T==`Tzero & phi1)
			 | (OP==`PHA & T==`Ttwo & phi1)
			 | (OP==`EOR_imm & T==`Tone & phi1)
			 | (OP==`EOR_imm & T==`Ttwo & phi1)
			 | (OP==`LSR & T==`Tone & phi1)
			 | (OP==`LSR & T==`Ttwo & phi1)
			 | (OP==`JMP_abs & T==`Ttwo & phi1)
			 | (OP==`EOR_abs & T==`Tzero & phi1)
			 | (OP==`EOR_abs & T==`Tone & phi1)
			 | (OP==`EOR_abs & T==`Ttwo & phi1)
			 | (OP==`LSR_abs & T==`Tzero & phi1)
			 | (OP==`LSR_abs & T==`Tone & phi1)
			 | (OP==`LSR_abs & T==`Ttwo & phi1)
			 | (OP==`LSR_abs & T==`Tfour & phi1)
			 | (OP==`LSR_abs & T==`Tfive & phi1)
			 | (OP==`BVC_rel & T==`Tzero & phi1)
			 | (OP==`BVC_rel & T==`Ttwo & phi1)
			 | (OP==`BVC_rel & T==`Tthree & phi1)
			 | (OP==`BVC_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BVC_rel & T==`T1BranchCross & phi1)
			 | (OP==`BVC_rel & T==`T1NoBranch & phi1)
			 | (OP==`EOR_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`EOR_izy & T==`Tone & phi1)
			 | (OP==`EOR_izy & T==`Ttwo & phi1)
			 | (OP==`EOR_izy & T==`Tfour & phi1)
			 | (OP==`EOR_zpx & T==`Tzero & phi1)
			 | (OP==`EOR_zpx & T==`Tone & phi1)
			 | (OP==`EOR_zpx & T==`Ttwo & phi1)
			 | (OP==`EOR_zpx & T==`Tthree & phi1)
			 | (OP==`LSR_zpx & T==`Tzero & phi1)
			 | (OP==`LSR_zpx & T==`Tone & phi1)
			 | (OP==`LSR_zpx & T==`Ttwo & phi1)
			 | (OP==`LSR_zpx & T==`Tthree & phi1)
			 | (OP==`LSR_zpx & T==`Tfour & phi1)
			 | (OP==`LSR_zpx & T==`Tfive & phi1)
			 | (OP==`CLI & T==`Tone & phi1)
			 | (OP==`CLI & T==`Ttwo & phi1)
			 | (OP==`EOR_aby & T==`TzeroNoCrossPg & phi1)
			 | (OP==`EOR_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`EOR_aby & T==`Tone & phi1)
			 | (OP==`EOR_aby & T==`Ttwo & phi1)
			 | (OP==`EOR_aby & T==`Tthree & phi1)
			 | (OP==`EOR_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`EOR_abx & T==`Tone & phi1)
			 | (OP==`EOR_abx & T==`Ttwo & phi1)
			 | (OP==`EOR_abx & T==`Tthree & phi1)
			 | (OP==`LSR_abx & T==`Tzero & phi1)
			 | (OP==`LSR_abx & T==`Tone & phi1)
			 | (OP==`LSR_abx & T==`Ttwo & phi1)
			 | (OP==`LSR_abx & T==`Tthree & phi1)
			 | (OP==`LSR_abx & T==`Tfive & phi1)
			 | (OP==`LSR_abx & T==`Tsix & phi1)
			 | (OP==`RTS & T==`Ttwo & phi1)
			 | (OP==`ADC_izx & T==`Tzero & phi1)
			 | (OP==`ADC_izx & T==`Tone & phi1)
			 | (OP==`ADC_izx & T==`Ttwo & phi1)
			 | (OP==`ADC_izx & T==`Tthree & phi1)
			 | (OP==`ADC_zp & T==`Tzero & phi1)
			 | (OP==`ADC_zp & T==`Tone & phi1)
			 | (OP==`ADC_zp & T==`Ttwo & phi1)
			 | (OP==`ROR_zp & T==`Tzero & phi1)
			 | (OP==`ROR_zp & T==`Tone & phi1)
			 | (OP==`ROR_zp & T==`Ttwo & phi1)
			 | (OP==`ROR_zp & T==`Tthree & phi1)
			 | (OP==`ROR_zp & T==`Tfour & phi1)
			 | (OP==`PLA & T==`Ttwo & phi1)
			 | (OP==`ADC_imm & T==`Tone & phi1)
			 | (OP==`ADC_imm & T==`Ttwo & phi1)
			 | (OP==`ROR & T==`Tone & phi1)
			 | (OP==`ROR & T==`Ttwo & phi1)
			 | (OP==`JMP_zp & T==`Ttwo & phi1)
			 | (OP==`ADC_abs & T==`Tzero & phi1)
			 | (OP==`ADC_abs & T==`Tone & phi1)
			 | (OP==`ADC_abs & T==`Ttwo & phi1)
			 | (OP==`ROR_abs & T==`Tzero & phi1)
			 | (OP==`ROR_abs & T==`Tone & phi1)
			 | (OP==`ROR_abs & T==`Ttwo & phi1)
			 | (OP==`ROR_abs & T==`Tfour & phi1)
			 | (OP==`ROR_abs & T==`Tfive & phi1)
			 | (OP==`BVS_rel & T==`Tzero & phi1)
			 | (OP==`BVS_rel & T==`Ttwo & phi1)
			 | (OP==`BVS_rel & T==`Tthree & phi1)
			 | (OP==`BVS_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BVS_rel & T==`T1BranchCross & phi1)
			 | (OP==`BVS_rel & T==`T1NoBranch & phi1)
			 | (OP==`ADC_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`ADC_izy & T==`Tone & phi1)
			 | (OP==`ADC_izy & T==`Ttwo & phi1)
			 | (OP==`ADC_izy & T==`Tfour & phi1)
			 | (OP==`ADC_zpx & T==`Tzero & phi1)
			 | (OP==`ADC_zpx & T==`Tone & phi1)
			 | (OP==`ADC_zpx & T==`Ttwo & phi1)
			 | (OP==`ADC_zpx & T==`Tthree & phi1)
			 | (OP==`ROR_zpx & T==`Tzero & phi1)
			 | (OP==`ROR_zpx & T==`Tone & phi1)
			 | (OP==`ROR_zpx & T==`Ttwo & phi1)
			 | (OP==`ROR_zpx & T==`Tthree & phi1)
			 | (OP==`ROR_zpx & T==`Tfour & phi1)
			 | (OP==`ROR_zpx & T==`Tfive & phi1)
			 | (OP==`SEI & T==`Tone & phi1)
			 | (OP==`SEI & T==`Ttwo & phi1)
			 | (OP==`ADC_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`ADC_aby & T==`Tone & phi1)
			 | (OP==`ADC_aby & T==`Ttwo & phi1)
			 | (OP==`ADC_aby & T==`Tthree & phi1)
			 | (OP==`ADC_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`ADC_abx & T==`Tone & phi1)
			 | (OP==`ADC_abx & T==`Ttwo & phi1)
			 | (OP==`ADC_abx & T==`Tthree & phi1)
			 | (OP==`ROR_abx & T==`Tzero & phi1)
			 | (OP==`ROR_abx & T==`Tone & phi1)
			 | (OP==`ROR_abx & T==`Ttwo & phi1)
			 | (OP==`ROR_abx & T==`Tthree & phi1)
			 | (OP==`ROR_abx & T==`Tfive & phi1)
			 | (OP==`ROR_abx & T==`Tsix & phi1)
			 | (OP==`STA_izx & T==`Tzero & phi1)
			 | (OP==`STA_izx & T==`Tone & phi1)
			 | (OP==`STA_izx & T==`Ttwo & phi1)
			 | (OP==`STA_izx & T==`Tthree & phi1)
			 | (OP==`STY_zp & T==`Tzero & phi1)
			 | (OP==`STY_zp & T==`Tone & phi1)
			 | (OP==`STY_zp & T==`Ttwo & phi1)
			 | (OP==`STA_zp & T==`Tzero & phi1)
			 | (OP==`STA_zp & T==`Tone & phi1)
			 | (OP==`STA_zp & T==`Ttwo & phi1)
			 | (OP==`STX_zp & T==`Tzero & phi1)
			 | (OP==`STX_zp & T==`Tone & phi1)
			 | (OP==`STX_zp & T==`Ttwo & phi1)
			 | (OP==`DEY & T==`Tone & phi1)
			 | (OP==`DEY & T==`Ttwo & phi1)
			 | (OP==`TXA & T==`Tone & phi1)
			 | (OP==`TXA & T==`Ttwo & phi1)
			 | (OP==`STY_abs & T==`Tzero & phi1)
			 | (OP==`STY_abs & T==`Tone & phi1)
			 | (OP==`STY_abs & T==`Ttwo & phi1)
			 | (OP==`STA_abs & T==`Tzero & phi1)
			 | (OP==`STA_abs & T==`Tone & phi1)
			 | (OP==`STA_abs & T==`Ttwo & phi1)
			 | (OP==`STX_abs & T==`Tzero & phi1)
			 | (OP==`STX_abs & T==`Tone & phi1)
			 | (OP==`STX_abs & T==`Ttwo & phi1)
			 | (OP==`BCC_rel & T==`Tzero & phi1)
			 | (OP==`BCC_rel & T==`Ttwo & phi1)
			 | (OP==`BCC_rel & T==`Tthree & phi1)
			 | (OP==`BCC_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BCC_rel & T==`T1BranchCross & phi1)
			 | (OP==`BCC_rel & T==`T1NoBranch & phi1)
			 | (OP==`STA_izy & T==`Tzero & phi1)
			 | (OP==`STA_izy & T==`Tone & phi1)
			 | (OP==`STA_izy & T==`Ttwo & phi1)
			 | (OP==`STA_izy & T==`Tfour & phi1)
			 | (OP==`STY_zpx & T==`Tzero & phi1)
			 | (OP==`STY_zpx & T==`Tone & phi1)
			 | (OP==`STY_zpx & T==`Ttwo & phi1)
			 | (OP==`STY_zpx & T==`Tthree & phi1)
			 | (OP==`STA_zpx & T==`Tzero & phi1)
			 | (OP==`STA_zpx & T==`Tone & phi1)
			 | (OP==`STA_zpx & T==`Ttwo & phi1)
			 | (OP==`STA_zpx & T==`Tthree & phi1)
			 | (OP==`STX_zpy & T==`Tzero & phi1)
			 | (OP==`STX_zpy & T==`Tone & phi1)
			 | (OP==`STX_zpy & T==`Ttwo & phi1)
			 | (OP==`STX_zpy & T==`Tthree & phi1)
			 | (OP==`TYA & T==`Tone & phi1)
			 | (OP==`TYA & T==`Ttwo & phi1)
			 | (OP==`STA_aby & T==`Tzero & phi1)
			 | (OP==`STA_aby & T==`Tone & phi1)
			 | (OP==`STA_aby & T==`Ttwo & phi1)
			 | (OP==`STA_aby & T==`Tthree & phi1)
			 | (OP==`TXS & T==`Tone & phi1)
			 | (OP==`TXS & T==`Ttwo & phi1)
			 | (OP==`STA_abx & T==`Tzero & phi1)
			 | (OP==`STA_abx & T==`Tone & phi1)
			 | (OP==`STA_abx & T==`Ttwo & phi1)
			 | (OP==`STA_abx & T==`Tthree & phi1)
			 | (OP==`LDY_imm & T==`Tone & phi1)
			 | (OP==`LDY_imm & T==`Ttwo & phi1)
			 | (OP==`LDA_izx & T==`Tzero & phi1)
			 | (OP==`LDA_izx & T==`Tone & phi1)
			 | (OP==`LDA_izx & T==`Ttwo & phi1)
			 | (OP==`LDA_izx & T==`Tthree & phi1)
			 | (OP==`LDX_imm & T==`Tone & phi1)
			 | (OP==`LDX_imm & T==`Ttwo & phi1)
			 | (OP==`LDY_zp & T==`Tzero & phi1)
			 | (OP==`LDY_zp & T==`Tone & phi1)
			 | (OP==`LDY_zp & T==`Ttwo & phi1)
			 | (OP==`LDA_zp & T==`Tzero & phi1)
			 | (OP==`LDA_zp & T==`Tone & phi1)
			 | (OP==`LDA_zp & T==`Ttwo & phi1)
			 | (OP==`LDX_zp & T==`Tzero & phi1)
			 | (OP==`LDX_zp & T==`Tone & phi1)
			 | (OP==`LDX_zp & T==`Ttwo & phi1)
			 | (OP==`TAY & T==`Tone & phi1)
			 | (OP==`TAY & T==`Ttwo & phi1)
			 | (OP==`LDA_imm & T==`Tone & phi1)
			 | (OP==`LDA_imm & T==`Ttwo & phi1)
			 | (OP==`TAX & T==`Tone & phi1)
			 | (OP==`TAX & T==`Ttwo & phi1)
			 | (OP==`LDY_abs & T==`Tzero & phi1)
			 | (OP==`LDY_abs & T==`Tone & phi1)
			 | (OP==`LDY_abs & T==`Ttwo & phi1)
			 | (OP==`LDA_abs & T==`Tzero & phi1)
			 | (OP==`LDA_abs & T==`Tone & phi1)
			 | (OP==`LDA_abs & T==`Ttwo & phi1)
			 | (OP==`LDX_abs & T==`Tzero & phi1)
			 | (OP==`LDX_abs & T==`Tone & phi1)
			 | (OP==`LDX_abs & T==`Ttwo & phi1)
			 | (OP==`BCS_rel & T==`Tzero & phi1)
			 | (OP==`BCS_rel & T==`Ttwo & phi1)
			 | (OP==`BCS_rel & T==`Tthree & phi1)
			 | (OP==`BCS_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BCS_rel & T==`T1BranchCross & phi1)
			 | (OP==`BCS_rel & T==`T1NoBranch & phi1)
			 | (OP==`LDA_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`LDA_izy & T==`Tone & phi1)
			 | (OP==`LDA_izy & T==`Ttwo & phi1)
			 | (OP==`LDA_izy & T==`Tfour & phi1)
			 | (OP==`LDY_zpx & T==`Tzero & phi1)
			 | (OP==`LDY_zpx & T==`Tone & phi1)
			 | (OP==`LDY_zpx & T==`Ttwo & phi1)
			 | (OP==`LDY_zpx & T==`Tthree & phi1)
			 | (OP==`LDA_zpx & T==`Tzero & phi1)
			 | (OP==`LDA_zpx & T==`Tone & phi1)
			 | (OP==`LDA_zpx & T==`Ttwo & phi1)
			 | (OP==`LDA_zpx & T==`Tthree & phi1)
			 | (OP==`LDX_zpy & T==`Tzero & phi1)
			 | (OP==`LDX_zpy & T==`Tone & phi1)
			 | (OP==`LDX_zpy & T==`Ttwo & phi1)
			 | (OP==`LDX_zpy & T==`Tthree & phi1)
			 | (OP==`CLV & T==`Tone & phi1)
			 | (OP==`CLV & T==`Ttwo & phi1)
			 | (OP==`LDA_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`LDA_aby & T==`Tone & phi1)
			 | (OP==`LDA_aby & T==`Ttwo & phi1)
			 | (OP==`LDA_aby & T==`Tthree & phi1)
			 | (OP==`TSX & T==`Tone & phi1)
			 | (OP==`TSX & T==`Ttwo & phi1)
			 | (OP==`LDY_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`LDY_abx & T==`Tone & phi1)
			 | (OP==`LDY_abx & T==`Ttwo & phi1)
			 | (OP==`LDY_abx & T==`Tthree & phi1)
			 | (OP==`LDA_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`LDA_abx & T==`Tone & phi1)
			 | (OP==`LDA_abx & T==`Ttwo & phi1)
			 | (OP==`LDA_abx & T==`Tthree & phi1)
			 | (OP==`LDX_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`LDX_aby & T==`Tone & phi1)
			 | (OP==`LDX_aby & T==`Ttwo & phi1)
			 | (OP==`LDX_aby & T==`Tthree & phi1)
			 | (OP==`CPY_imm & T==`Tone & phi1)
			 | (OP==`CPY_imm & T==`Ttwo & phi1)
			 | (OP==`CMP_izx & T==`Tzero & phi1)
			 | (OP==`CMP_izx & T==`Tone & phi1)
			 | (OP==`CMP_izx & T==`Ttwo & phi1)
			 | (OP==`CMP_izx & T==`Tthree & phi1)
			 | (OP==`CPY_zp & T==`Tzero & phi1)
			 | (OP==`CPY_zp & T==`Tone & phi1)
			 | (OP==`CPY_zp & T==`Ttwo & phi1)
			 | (OP==`CMP_zp & T==`Tzero & phi1)
			 | (OP==`CMP_zp & T==`Tone & phi1)
			 | (OP==`CMP_zp & T==`Ttwo & phi1)
			 | (OP==`DEC_zp & T==`Tzero & phi1)
			 | (OP==`DEC_zp & T==`Tone & phi1)
			 | (OP==`DEC_zp & T==`Ttwo & phi1)
			 | (OP==`DEC_zp & T==`Tthree & phi1)
			 | (OP==`DEC_zp & T==`Tfour & phi1)
			 | (OP==`INY & T==`Tone & phi1)
			 | (OP==`INY & T==`Ttwo & phi1)
			 | (OP==`CMP_imm & T==`Tone & phi1)
			 | (OP==`CMP_imm & T==`Ttwo & phi1)
			 | (OP==`DEX & T==`Tone & phi1)
			 | (OP==`DEX & T==`Ttwo & phi1)
			 | (OP==`CPY_abs & T==`Tzero & phi1)
			 | (OP==`CPY_abs & T==`Tone & phi1)
			 | (OP==`CPY_abs & T==`Ttwo & phi1)
			 | (OP==`CMP_abs & T==`Tzero & phi1)
			 | (OP==`CMP_abs & T==`Tone & phi1)
			 | (OP==`CMP_abs & T==`Ttwo & phi1)
			 | (OP==`DEC_abs & T==`Tzero & phi1)
			 | (OP==`DEC_abs & T==`Tone & phi1)
			 | (OP==`DEC_abs & T==`Ttwo & phi1)
			 | (OP==`DEC_abs & T==`Tfour & phi1)
			 | (OP==`DEC_abs & T==`Tfive & phi1)
			 | (OP==`BNE_rel & T==`Tzero & phi1)
			 | (OP==`BNE_rel & T==`Ttwo & phi1)
			 | (OP==`BNE_rel & T==`Tthree & phi1)
			 | (OP==`BNE_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BNE_rel & T==`T1BranchCross & phi1)
			 | (OP==`BNE_rel & T==`T1NoBranch & phi1)
			 | (OP==`CMP_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`CMP_izy & T==`Tone & phi1)
			 | (OP==`CMP_izy & T==`Ttwo & phi1)
			 | (OP==`CMP_izy & T==`Tfour & phi1)
			 | (OP==`CMP_zpx & T==`Tzero & phi1)
			 | (OP==`CMP_zpx & T==`Tone & phi1)
			 | (OP==`CMP_zpx & T==`Ttwo & phi1)
			 | (OP==`CMP_zpx & T==`Tthree & phi1)
			 | (OP==`DEC_zpx & T==`Tzero & phi1)
			 | (OP==`DEC_zpx & T==`Tone & phi1)
			 | (OP==`DEC_zpx & T==`Ttwo & phi1)
			 | (OP==`DEC_zpx & T==`Tthree & phi1)
			 | (OP==`DEC_zpx & T==`Tfour & phi1)
			 | (OP==`DEC_zpx & T==`Tfive & phi1)
			 | (OP==`CLD & T==`Tone & phi1)
			 | (OP==`CLD & T==`Ttwo & phi1)
			 | (OP==`CMP_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`CMP_aby & T==`Tone & phi1)
			 | (OP==`CMP_aby & T==`Ttwo & phi1)
			 | (OP==`CMP_aby & T==`Tthree & phi1)
			 | (OP==`CMP_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`CMP_abx & T==`Tone & phi1)
			 | (OP==`CMP_abx & T==`Ttwo & phi1)
			 | (OP==`CMP_abx & T==`Tthree & phi1)
			 | (OP==`DEC_abx & T==`Tzero & phi1)
			 | (OP==`DEC_abx & T==`Tone & phi1)
			 | (OP==`DEC_abx & T==`Ttwo & phi1)
			 | (OP==`DEC_abx & T==`Tthree & phi1)
			 | (OP==`DEC_abx & T==`Tfive & phi1)
			 | (OP==`DEC_abx & T==`Tsix & phi1)
			 | (OP==`CPX_imm & T==`Tone & phi1)
			 | (OP==`CPX_imm & T==`Ttwo & phi1)
			 | (OP==`SBC_izx & T==`Tzero & phi1)
			 | (OP==`SBC_izx & T==`Tone & phi1)
			 | (OP==`SBC_izx & T==`Ttwo & phi1)
			 | (OP==`SBC_izx & T==`Tthree & phi1)
			 | (OP==`CPX_zp & T==`Tzero & phi1)
			 | (OP==`CPX_zp & T==`Tone & phi1)
			 | (OP==`CPX_zp & T==`Ttwo & phi1)
			 | (OP==`SBC_zp & T==`Tzero & phi1)
			 | (OP==`SBC_zp & T==`Tone & phi1)
			 | (OP==`SBC_zp & T==`Ttwo & phi1)
			 | (OP==`INC_zp & T==`Tzero & phi1)
			 | (OP==`INC_zp & T==`Tone & phi1)
			 | (OP==`INC_zp & T==`Ttwo & phi1)
			 | (OP==`INC_zp & T==`Tthree & phi1)
			 | (OP==`INX & T==`Tone & phi1)
			 | (OP==`INX & T==`Ttwo & phi1)
			 | (OP==`SBC_imm & T==`Tone & phi1)
			 | (OP==`SBC_imm & T==`Ttwo & phi1)
			 | (OP==`NOP & T==`Tone & phi1)
			 | (OP==`NOP & T==`Ttwo & phi1)
			 | (OP==`CPX_abs & T==`Tzero & phi1)
			 | (OP==`CPX_abs & T==`Tone & phi1)
			 | (OP==`CPX_abs & T==`Ttwo & phi1)
			 | (OP==`SBC_abs & T==`Tzero & phi1)
			 | (OP==`SBC_abs & T==`Tone & phi1)
			 | (OP==`SBC_abs & T==`Ttwo & phi1)
			 | (OP==`INC_abs & T==`Tzero & phi1)
			 | (OP==`INC_abs & T==`Tone & phi1)
			 | (OP==`INC_abs & T==`Ttwo & phi1)
			 | (OP==`INC_abs & T==`Tfour & phi1)
			 | (OP==`BEQ_rel & T==`Tzero & phi1)
			 | (OP==`BEQ_rel & T==`Ttwo & phi1)
			 | (OP==`BEQ_rel & T==`Tthree & phi1)
			 | (OP==`BEQ_rel & T==`T1BranchNoCross & phi1)
			 | (OP==`BEQ_rel & T==`T1BranchCross & phi1)
			 | (OP==`BEQ_rel & T==`T1NoBranch & phi1)
			 | (OP==`SBC_izy & T==`TzeroCrossPg & phi1)
			 | (OP==`SBC_izy & T==`Tone & phi1)
			 | (OP==`SBC_izy & T==`Ttwo & phi1)
			 | (OP==`SBC_izy & T==`Tfour & phi1)
			 | (OP==`SBC_zpx & T==`Tzero & phi1)
			 | (OP==`SBC_zpx & T==`Tone & phi1)
			 | (OP==`SBC_zpx & T==`Ttwo & phi1)
			 | (OP==`SBC_zpx & T==`Tthree & phi1)
			 | (OP==`INC_zpx & T==`Tzero & phi1)
			 | (OP==`INC_zpx & T==`Tone & phi1)
			 | (OP==`INC_zpx & T==`Ttwo & phi1)
			 | (OP==`INC_zpx & T==`Tthree & phi1)
			 | (OP==`INC_zpx & T==`Tfour & phi1)
			 | (OP==`SED & T==`Tone & phi1)
			 | (OP==`SED & T==`Ttwo & phi1)
			 | (OP==`SBC_aby & T==`TzeroCrossPg & phi1)
			 | (OP==`SBC_aby & T==`Tone & phi1)
			 | (OP==`SBC_aby & T==`Ttwo & phi1)
			 | (OP==`SBC_aby & T==`Tthree & phi1)
			 | (OP==`SBC_abx & T==`TzeroCrossPg & phi1)
			 | (OP==`SBC_abx & T==`Tone & phi1)
			 | (OP==`SBC_abx & T==`Ttwo & phi1)
			 | (OP==`SBC_abx & T==`Tthree & phi1)
			 | (OP==`INC_abx & T==`Tzero & phi1)
			 | (OP==`INC_abx & T==`Tone & phi1)
			 | (OP==`INC_abx & T==`Ttwo & phi1)
			 | (OP==`INC_abx & T==`Tthree & phi1)
			 | (OP==`INC_abx & T==`Tfive & phi1)
			;

    assign control[`SB_AC] = (OP==`PLA & T==`Tone & phi1)
         | (OP==`TXA & T==`Tone & phi1)
         | (OP==`TYA & T==`Tone & phi1)
         | (OP==`LDA_izx & T==`Tone & phi1)
         | (OP==`LDA_zp & T==`Tone & phi1)
         | (OP==`LDA_imm & T==`Tone & phi1)
         | (OP==`LDA_abs & T==`Tone & phi1)
         | (OP==`LDA_izy & T==`Tone & phi1)
         | (OP==`LDA_zpx & T==`Tone & phi1)
         | (OP==`LDA_aby & T==`Tone & phi1)
         | (OP==`LDA_abx & T==`Tone & phi1)
         | ((T==`Ttwo) & (prevOP == `ADC_abs || prevOP == `ADC_abx || prevOP == `ADC_aby || prevOP == `ADC_imm || 
             prevOP == `ADC_izx || prevOP == `ADC_izy || prevOP == `ADC_zp  || prevOP == `ADC_zpx ||
             prevOP == `SBC_abs || prevOP == `SBC_abx || prevOP == `SBC_aby || prevOP == `SBC_imm || 
             prevOP == `SBC_izx || prevOP == `SBC_izy || prevOP == `SBC_zp  || prevOP == `SBC_zpx ||
             prevOP == `AND_imm || prevOP == `AND_abs || prevOP == `AND_abx || prevOP == `AND_aby ||
             prevOP == `AND_izx || prevOP == `AND_izy || prevOP == `AND_zp  || prevOP == `AND_zpx ||
             prevOP == `ORA_imm || prevOP == `ORA_abs || prevOP == `ORA_abx || prevOP == `ORA_aby ||
             prevOP == `ORA_izx || prevOP == `ORA_izy || prevOP == `ORA_zp  || prevOP == `ORA_zpx ||
             prevOP == `EOR_imm || prevOP == `EOR_abs || prevOP == `EOR_abx || prevOP == `EOR_aby ||
             prevOP == `EOR_izx || prevOP == `EOR_izy || prevOP == `EOR_zp  || prevOP == `EOR_zpx ||
             prevOP == `ASL     || prevOP == `LSR     || prevOP == `ROL     || prevOP == `ROR     ))
                ;

assign control[`AC_DB] = (OP==`PHA & T==`Tzero & phi1)
			 | (OP==`STA_izx & T==`Tzero & phi1)
			 | (OP==`STA_zp & T==`Tzero & phi1)
			 | (OP==`STA_abs & T==`Tzero & phi1)
			 | (OP==`STA_izy & T==`Tzero & phi1)
			 | (OP==`STA_zpx & T==`Tzero & phi1)
			 | (OP==`STA_aby & T==`Tzero & phi1)
			 | (OP==`STA_abx & T==`Tzero & phi1)
			;

assign control[`AC_SB] = (OP==`ORA_izx & T==`Tone & phi1)
			 | (OP==`ORA_zp & T==`Tone & phi1)
			 | (OP==`ORA_imm & T==`Tone & phi1)
			 | (OP==`ASL & T==`Tone & phi1)
			 | (OP==`ORA_abs & T==`Tone & phi1)
			 | (OP==`ORA_izy & T==`Tone & phi1)
			 | (OP==`ORA_zpx & T==`Tone & phi1)
			 | (OP==`ORA_aby & T==`Tone & phi1)
			 | (OP==`ORA_abx & T==`Tone & phi1)
			 | (OP==`AND_izx & T==`Tone & phi1)
			 | (OP==`BIT_zp & T==`Tone & phi1)
			 | (OP==`AND_zp & T==`Tone & phi1)
			 | (OP==`AND_imm & T==`Tone & phi1)
			 | (OP==`ROL & T==`Tone & phi1)
			 | (OP==`BIT_abs & T==`Tone & phi1)
			 | (OP==`AND_abs & T==`Tone & phi1)
			 | (OP==`AND_izy & T==`Tone & phi1)
			 | (OP==`AND_zpx & T==`Tone & phi1)
			 | (OP==`AND_aby & T==`Tone & phi1)
			 | (OP==`AND_abx & T==`Tone & phi1)
			 | (OP==`EOR_izx & T==`Tone & phi1)
			 | (OP==`EOR_zp & T==`Tone & phi1)
			 | (OP==`EOR_imm & T==`Tone & phi1)
			 | (OP==`LSR & T==`Tone & phi1)
			 | (OP==`EOR_abs & T==`Tone & phi1)
			 | (OP==`EOR_izy & T==`Tone & phi1)
			 | (OP==`EOR_zpx & T==`Tone & phi1)
			 | (OP==`EOR_aby & T==`Tone & phi1)
			 | (OP==`EOR_abx & T==`Tone & phi1)
			 | (OP==`ADC_izx & T==`Tone & phi1)
			 | (OP==`ADC_zp & T==`Tone & phi1)
			 | (OP==`ADC_imm & T==`Tone & phi1)
			 | (OP==`ROR & T==`Tone & phi1)
			 | (OP==`ADC_abs & T==`Tone & phi1)
			 | (OP==`ADC_izy & T==`Tone & phi1)
			 | (OP==`ADC_zpx & T==`Tone & phi1)
			 | (OP==`ADC_aby & T==`Tone & phi1)
			 | (OP==`ADC_abx & T==`Tone & phi1)
			 | (OP==`STA_izx & T==`Tone & phi1)
			 | (OP==`STA_zp & T==`Tone & phi1)
			 | (OP==`STA_abs & T==`Tone & phi1)
			 | (OP==`STA_izy & T==`Tone & phi1)
			 | (OP==`STA_zpx & T==`Tone & phi1)
			 | (OP==`STA_aby & T==`Tone & phi1)
			 | (OP==`STA_abx & T==`Tone & phi1)
			 | (OP==`TAY & T==`Tone & phi1)
			 | (OP==`TAX & T==`Tone & phi1)
			 | (OP==`CMP_izx & T==`Tone & phi1)
			 | (OP==`CMP_zp & T==`Tone & phi1)
			 | (OP==`CMP_imm & T==`Tone & phi1)
			 | (OP==`CMP_abs & T==`Tone & phi1)
			 | (OP==`CMP_izy & T==`Tone & phi1)
			 | (OP==`CMP_zpx & T==`Tone & phi1)
			 | (OP==`CMP_aby & T==`Tone & phi1)
			 | (OP==`CMP_abx & T==`Tone & phi1)
			 | (OP==`SBC_izx & T==`Tone & phi1)
			 | (OP==`SBC_zp & T==`Tone & phi1)
			 | (OP==`SBC_imm & T==`Tone & phi1)
			 | (OP==`SBC_abs & T==`Tone & phi1)
			 | (OP==`SBC_izy & T==`Tone & phi1)
			 | (OP==`SBC_zpx & T==`Tone & phi1)
			 | (OP==`SBC_aby & T==`Tone & phi1)
			 | (OP==`SBC_abx & T==`Tone & phi1)
			;

    assign control[`SB_X] = (OP==`LDX_imm & T==`Tone & phi1)
                 | (OP==`LDX_zp & T==`Tone & phi1)
                 | (OP==`TAX & T==`Tone & phi1)
                 | (OP==`LDX_abs & T==`Tone & phi1)
                 | (OP==`LDX_zpy & T==`Tone & phi1)
                 | (OP==`TSX & T==`Tone & phi1)
                 | (OP==`LDX_aby & T==`Tone & phi1)
                 | ((T==`Ttwo) & (prevOP == `INX || prevOP == `DEX))
                ;

assign control[`X_SB] = (OP==`ORA_izx & T==`Tthree & phi1)
			 | (OP==`ORA_zpx & T==`Tthree & phi1)
			 | (OP==`ASL_zpx & T==`Tthree & phi1)
			 | (OP==`ORA_abx & T==`Tthree & phi1)
			 | (OP==`ASL_abx & T==`Tthree & phi1)
			 | (OP==`AND_izx & T==`Tthree & phi1)
			 | (OP==`AND_zpx & T==`Tthree & phi1)
			 | (OP==`ROL_zpx & T==`Tthree & phi1)
			 | (OP==`AND_abx & T==`Tthree & phi1)
			 | (OP==`ROL_abx & T==`Tthree & phi1)
			 | (OP==`EOR_izx & T==`Tthree & phi1)
			 | (OP==`EOR_zpx & T==`Tthree & phi1)
			 | (OP==`LSR_zpx & T==`Tthree & phi1)
			 | (OP==`EOR_abx & T==`Tthree & phi1)
			 | (OP==`LSR_abx & T==`Tthree & phi1)
			 | (OP==`ADC_izx & T==`Tthree & phi1)
			 | (OP==`ADC_zpx & T==`Tthree & phi1)
			 | (OP==`ROR_zpx & T==`Tthree & phi1)
			 | (OP==`ADC_abx & T==`Tthree & phi1)
			 | (OP==`ROR_abx & T==`Tthree & phi1)
			 | (OP==`STA_izx & T==`Tthree & phi1)
			 | (OP==`STX_zp & T==`Tzero & phi1)
			 | (OP==`TXA & T==`Tone & phi1)
			 | (OP==`STX_abs & T==`Tzero & phi1)
			 | (OP==`STY_zpx & T==`Tthree & phi1)
			 | (OP==`STA_zpx & T==`Tthree & phi1)
			 | (OP==`STX_zpy & T==`Tzero & phi1)
			 | (OP==`TXS & T==`Tone & phi1)
			 | (OP==`STA_abx & T==`Tthree & phi1)
			 | (OP==`LDA_izx & T==`Tthree & phi1)
			 | (OP==`LDY_zpx & T==`Tthree & phi1)
			 | (OP==`LDA_zpx & T==`Tthree & phi1)
			 | (OP==`LDY_abx & T==`Tthree & phi1)
			 | (OP==`LDA_abx & T==`Tthree & phi1)
			 | (OP==`CMP_izx & T==`Tthree & phi1)
			 | (OP==`DEX & T==`Tone & phi1)
			 | (OP==`CMP_zpx & T==`Tthree & phi1)
			 | (OP==`DEC_zpx & T==`Tthree & phi1)
			 | (OP==`CMP_abx & T==`Tthree & phi1)
			 | (OP==`DEC_abx & T==`Tthree & phi1)
			 | (OP==`CPX_imm & T==`Tone & phi1)
			 | (OP==`SBC_izx & T==`Tthree & phi1)
			 | (OP==`CPX_zp & T==`Tone & phi1)
			 | (OP==`INX & T==`Tone & phi1)
			 | (OP==`CPX_abs & T==`Tone & phi1)
			 | (OP==`SBC_zpx & T==`Tthree & phi1)
			 | (OP==`INC_zpx & T==`Tthree & phi1)
			 | (OP==`SBC_abx & T==`Tthree & phi1)
			 | (OP==`INC_abx & T==`Tthree & phi1)
			;

    assign control[`SB_Y] = (OP==`LDY_imm & T==`Tone & phi1)
                 | (OP==`LDY_zp & T==`Tone & phi1)
                 | (OP==`TAY & T==`Tone & phi1)
                 | (OP==`LDY_abs & T==`Tone & phi1)
                 | (OP==`LDY_zpx & T==`Tone & phi1)
                 | (OP==`LDY_abx & T==`Tone & phi1)
                 | ((T==`Ttwo) & (prevOP == `INY || prevOP == `DEY))
                ;  

assign control[`Y_SB] = (OP==`ORA_izy & T==`Tfour & phi1)
			 | (OP==`ORA_aby & T==`Tthree & phi1)
			 | (OP==`AND_izy & T==`Tfour & phi1)
			 | (OP==`AND_aby & T==`Tthree & phi1)
			 | (OP==`EOR_izy & T==`Tfour & phi1)
			 | (OP==`EOR_aby & T==`Tthree & phi1)
			 | (OP==`ADC_izy & T==`Tfour & phi1)
			 | (OP==`ADC_aby & T==`Tthree & phi1)
			 | (OP==`STY_zp & T==`Tzero & phi1)
			 | (OP==`DEY & T==`Tone & phi1)
			 | (OP==`STY_abs & T==`Tzero & phi1)
			 | (OP==`STA_izy & T==`Tfour & phi1)
			 | (OP==`STY_zpx & T==`Tzero & phi1)
			 | (OP==`STX_zpy & T==`Tthree & phi1)
			 | (OP==`TYA & T==`Tone & phi1)
			 | (OP==`STA_aby & T==`Tthree & phi1)
			 | (OP==`LDA_izy & T==`Tfour & phi1)
			 | (OP==`LDX_zpy & T==`Tthree & phi1)
			 | (OP==`LDA_aby & T==`Tthree & phi1)
			 | (OP==`LDX_aby & T==`Tthree & phi1)
			 | (OP==`CPY_imm & T==`Tone & phi1)
			 | (OP==`CPY_zp & T==`Tone & phi1)
			 | (OP==`INY & T==`Tone & phi1)
			 | (OP==`CPY_abs & T==`Tone & phi1)
			 | (OP==`CMP_izy & T==`Tfour & phi1)
			 | (OP==`CMP_aby & T==`Tthree & phi1)
			 | (OP==`SBC_izy & T==`Tfour & phi1)
			 | (OP==`SBC_aby & T==`Tthree & phi1)
			;

assign control[`P_DB] = (OP==`BRK & T==`Tfour & phi2)
			 | (OP==`BRK & T==`Tfive & phi1)
			 | (OP==`PHP & T==`Tzero & phi1)
			 | (OP==`PHP & T==`Ttwo & phi2)
			;

assign control[`DB_P] = (OP==`PLP & T==`Tzero & phi2)
			 | (OP==`PLP & T==`Tone & phi1)
			 | (OP==`RTI & T==`Tfour & phi2)
			 | (OP==`RTI & T==`Tfive & phi1)
			;

assign control[`SET_C] = (OP==`SEC & T==`Tone & phi1)
			 | (OP==`SEC & T==`Ttwo & phi2)
			;

assign control[`CLR_C] = (OP==`CLC & T==`Tone & phi1)
			 | (OP==`CLC & T==`Ttwo & phi2)
			;

assign control[`SET_I] = (OP==`BRK & T==`Tzero)
			 | (OP==`SEI & T==`Tone & phi1)
			 | (OP==`SEI & T==`Ttwo & phi2)
			;

assign control[`CLR_I] = (OP==`CLI & T==`Tone & phi1)
			 | (OP==`CLI & T==`Ttwo & phi2)
			;

assign control[`CLR_V] = (OP==`CLV & T==`Tone & phi1)
			 | (OP==`CLV & T==`Ttwo & phi2)
			;

assign control[`SET_D] = (OP==`SED & T==`Tone & phi1)
			 | (OP==`SED & T==`Ttwo & phi2)
			;

assign control[`CLR_D] = (OP==`CLD & T==`Tone & phi1)
			 | (OP==`CLD & T==`Ttwo & phi2)
			;


assign control[`FLAG_DBZ] = (OP==`BIT_zp & T==`Tone & phi2)
			;

assign control[`FLAG_DB] = (OP==`BIT_zp & T==`Tzero & phi2)
			 | (OP==`DEY & T==`Tone & phi2)
			 | (OP==`TXA & T==`Tone & phi1)
			 | (OP==`TYA & T==`Tone & phi1)
			 | (OP==`TXS & T==`Tone & phi1)
			 | (OP==`LDY_imm & T==`Ttwo & phi2)
			 | (OP==`LDA_izx & T==`Tzero & phi2)
			 | (OP==`LDX_imm & T==`Ttwo & phi2)
			 | (OP==`LDY_zp & T==`Tzero & phi2)
			 | (OP==`LDA_zp & T==`Tzero & phi2)
			 | (OP==`LDX_zp & T==`Tzero & phi2)
			 | (OP==`TAY & T==`Tone & phi1)
			 | (OP==`LDA_imm & T==`Ttwo & phi2)
			 | (OP==`TAX & T==`Tone & phi1)
			 | (OP==`LDY_abs & T==`Tzero & phi2)
			 | (OP==`LDA_abs & T==`Tzero & phi2)
			 | (OP==`LDX_abs & T==`Tzero & phi2)
			 | (OP==`LDA_izy & T==`TzeroNoCrossPg & phi2)
			 | (OP==`LDA_izy & T==`TzeroCrossPg & phi2)
			 | (OP==`LDY_zpx & T==`Tzero & phi2)
			 | (OP==`LDA_zpx & T==`Tzero & phi2)
			 | (OP==`LDX_zpy & T==`Tzero & phi2)
			 | (OP==`LDA_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`LDA_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`TSX & T==`Tone & phi1)
			 | (OP==`LDY_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`LDY_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`LDA_abx & T==`TzeroNoCrossPg & phi2)
			 | (OP==`LDA_abx & T==`TzeroCrossPg & phi2)
			 | (OP==`LDX_aby & T==`TzeroNoCrossPg & phi2)
			 | (OP==`LDX_aby & T==`TzeroCrossPg & phi2)
			 | (OP==`DEC_zp & T==`Tfour & phi2)
			 | (OP==`INY & T==`Tone & phi2)
			 | (OP==`DEX & T==`Tone & phi2)
			 | (OP==`DEC_abs & T==`Tfive & phi2)
			 | (OP==`DEC_zpx & T==`Tfive & phi2)
			 | (OP==`DEC_abx & T==`Tsix & phi2)
			 | (OP==`INC_zp & T==`Tfour & phi2)
			 | (OP==`INX & T==`Tone & phi2)
			 | (OP==`INC_abs & T==`Tfive & phi2)
			 | (OP==`INC_zpx & T==`Tfive & phi2)
			 | (OP==`INC_abx & T==`Tsix & phi2)
			;

assign control[`FLAG_ALU] = (OP==`ORA_izx & T==`Tone & phi2)
			 | (OP==`ORA_zp & T==`Tone & phi2)
			 | (OP==`ASL_zp & T==`Tfour & phi2)
			 | (OP==`ORA_imm & T==`Tone & phi2)
			 | (OP==`ASL & T==`Tone & phi2)
			 | (OP==`ORA_abs & T==`Tone & phi2)
			 | (OP==`ASL_abs & T==`Tfive & phi2)
			 | (OP==`ORA_izy & T==`Tone & phi2)
			 | (OP==`ORA_zpx & T==`Tone & phi2)
			 | (OP==`ASL_zpx & T==`Tfive & phi2)
			 | (OP==`ORA_aby & T==`Tone & phi2)
			 | (OP==`ORA_abx & T==`Tone & phi2)
			 | (OP==`ASL_abx & T==`Tsix & phi2)
			 | (OP==`AND_izx & T==`Tone & phi2)
			 | (OP==`AND_zp & T==`Tone & phi2)
			 | (OP==`ROL_zp & T==`Tfour & phi2)
			 | (OP==`AND_imm & T==`Tone & phi2)
			 | (OP==`ROL & T==`Tone & phi2)
			 | (OP==`AND_abs & T==`Tone & phi2)
			 | (OP==`ROL_abs & T==`Tfive & phi2)
			 | (OP==`AND_izy & T==`Tone & phi2)
			 | (OP==`AND_zpx & T==`Tone & phi2)
			 | (OP==`ROL_zpx & T==`Tfive & phi2)
			 | (OP==`AND_aby & T==`Tone & phi2)
			 | (OP==`AND_abx & T==`Tone & phi2)
			 | (OP==`ROL_abx & T==`Tsix & phi2)
			 | (OP==`EOR_izx & T==`Tone & phi2)
			 | (OP==`EOR_zp & T==`Tone & phi2)
			 | (OP==`LSR_zp & T==`Tone & phi2)
			 | (OP==`LSR_zp & T==`Tfour & phi2)
			 | (OP==`EOR_imm & T==`Tone & phi2)
			 | (OP==`LSR & T==`Tone & phi2)
			 | (OP==`EOR_abs & T==`Tone & phi2)
			 | (OP==`LSR_abs & T==`Tone & phi2)
			 | (OP==`LSR_abs & T==`Tfive & phi2)
			 | (OP==`EOR_izy & T==`Tone & phi2)
			 | (OP==`EOR_zpx & T==`Tone & phi2)
			 | (OP==`LSR_zpx & T==`Tone & phi2)
			 | (OP==`LSR_zpx & T==`Tfive & phi2)
			 | (OP==`EOR_aby & T==`Tone & phi2)
			 | (OP==`EOR_abx & T==`Tone & phi2)
			 | (OP==`LSR_abx & T==`Tone & phi2)
			 | (OP==`LSR_abx & T==`Tsix & phi2)
			 | (OP==`ADC_izx & T==`Tone & phi2)
			 | (OP==`ADC_zp & T==`Tone & phi2)
			 | (OP==`ROR_zp & T==`Tfour & phi2)
			 | (OP==`ADC_imm & T==`Tone & phi2)
			 | (OP==`ROR & T==`Tone & phi2)
			 | (OP==`ADC_abs & T==`Tone & phi2)
			 | (OP==`ROR_abs & T==`Tfive & phi2)
			 | (OP==`ADC_izy & T==`Tone & phi2)
			 | (OP==`ADC_zpx & T==`Tone & phi2)
			 | (OP==`ROR_zpx & T==`Tfive & phi2)
			 | (OP==`ADC_aby & T==`Tone & phi2)
			 | (OP==`ADC_abx & T==`Tone & phi2)
			 | (OP==`ROR_abx & T==`Tsix & phi2)
			 | (OP==`CPY_imm & T==`Tone & phi2)
			 | (OP==`CMP_izx & T==`Tone & phi2)
			 | (OP==`CPY_zp & T==`Tone & phi2)
			 | (OP==`CMP_zp & T==`Tone & phi2)
			 | (OP==`CMP_imm & T==`Tone & phi2)
			 | (OP==`CPY_abs & T==`Tone & phi2)
			 | (OP==`CMP_abs & T==`Tone & phi2)
			 | (OP==`CMP_izy & T==`Tone & phi2)
			 | (OP==`CMP_zpx & T==`Tone & phi2)
			 | (OP==`CMP_aby & T==`Tone & phi2)
			 | (OP==`CMP_abx & T==`Tone & phi2)
			 | (OP==`CPX_imm & T==`Tone & phi2)
			 | (OP==`SBC_izx & T==`Tone & phi2)
			 | (OP==`CPX_zp & T==`Tone & phi2)
			 | (OP==`SBC_zp & T==`Tone & phi2)
			 | (OP==`SBC_imm & T==`Tone & phi2)
			 | (OP==`CPX_abs & T==`Tone & phi2)
			 | (OP==`SBC_abs & T==`Tone & phi2)
			 | (OP==`SBC_izy & T==`Tone & phi2)
			 | (OP==`SBC_zpx & T==`Tone & phi2)
			 | (OP==`SBC_aby & T==`Tone & phi2)
			 | (OP==`SBC_abx & T==`Tone & phi2)
			;

assign control[`nRW] = (OP==`BRK & T==`Tthree & activeInt != `RST_i)
			|(OP==`BRK & T==`Tfour & activeInt != `RST_i)
			|(OP==`BRK & T==`Tfive & activeInt != `RST_i)
			 | (OP==`ASL_zp & T==`Tzero)
			 | (OP==`ASL_zp & T==`Tfour)
			 | (OP==`PHP & T==`Tzero)
			 | (OP==`ASL_abs & T==`Tzero)
			 | (OP==`ASL_abs & T==`Tfive)
			 | (OP==`ASL_zpx & T==`Tzero)
			 | (OP==`ASL_zpx & T==`Tfive)
			 | (OP==`ASL_abx & T==`Tzero)
			 | (OP==`ASL_abx & T==`Tsix)
			 | (OP==`JSR_abs & T==`Tfour)
			 | (OP==`JSR_abs & T==`Tfive)
			 | (OP==`ROL_zp & T==`Tzero)
			 | (OP==`ROL_zp & T==`Tfour)
			 | (OP==`ROL_abs & T==`Tzero)
			 | (OP==`ROL_abs & T==`Tfive)
			 | (OP==`ROL_zpx & T==`Tzero)
			 | (OP==`ROL_zpx & T==`Tfive)
			 | (OP==`ROL_abx & T==`Tzero)
			 | (OP==`ROL_abx & T==`Tsix)
			 | (OP==`LSR_zp & T==`Tzero)
			 | (OP==`LSR_zp & T==`Tfour)
			 | (OP==`PHA & T==`Tzero)
			 | (OP==`LSR_abs & T==`Tzero)
			 | (OP==`LSR_abs & T==`Tfive)
			 | (OP==`LSR_zpx & T==`Tzero)
			 | (OP==`LSR_zpx & T==`Tfive)
			 | (OP==`LSR_abx & T==`Tzero)
			 | (OP==`LSR_abx & T==`Tsix)
			 | (OP==`ROR_zp & T==`Tzero)
			 | (OP==`ROR_zp & T==`Tfour)
			 | (OP==`ROR_abs & T==`Tzero)
			 | (OP==`ROR_abs & T==`Tfive)
			 | (OP==`ROR_zpx & T==`Tzero)
			 | (OP==`ROR_zpx & T==`Tfive)
			 | (OP==`ROR_abx & T==`Tzero)
			 | (OP==`ROR_abx & T==`Tsix)
			 | (OP==`STA_izx & T==`Tzero)
			 | (OP==`STY_zp & T==`Tzero)
			 | (OP==`STA_zp & T==`Tzero)
			 | (OP==`STX_zp & T==`Tzero)
			 | (OP==`STY_abs & T==`Tzero)
			 | (OP==`STA_abs & T==`Tzero)
			 | (OP==`STX_abs & T==`Tzero)
			 | (OP==`STA_izy & T==`Tzero)
			 | (OP==`STY_zpx & T==`Tzero)
			 | (OP==`STA_zpx & T==`Tzero)
			 | (OP==`STX_zpy & T==`Tzero)
			 | (OP==`STA_aby & T==`Tzero)
			 | (OP==`STA_abx & T==`Tzero)
			 | (OP==`DEC_zp & T==`Tzero)
			 | (OP==`DEC_zp & T==`Tfour)
			 | (OP==`DEC_abs & T==`Tzero)
			 | (OP==`DEC_abs & T==`Tfive)
			 | (OP==`DEC_zpx & T==`Tzero)
			 | (OP==`DEC_zpx & T==`Tfive)
			 | (OP==`DEC_abx & T==`Tzero)
			 | (OP==`DEC_abx & T==`Tsix)
			 | (OP==`INC_zp & T==`Tzero)
			 | (OP==`INC_zp & T==`Tfour)
			 | (OP==`INC_abs & T==`Tzero)
			 | (OP==`INC_abs & T==`Tfive)
			 | (OP==`INC_zpx & T==`Tzero)
			 | (OP==`INC_zpx & T==`Tfive)
			 | (OP==`INC_abx & T==`Tzero)
			 | (OP==`INC_abx & T==`Tsix)
			;
 
endmodule