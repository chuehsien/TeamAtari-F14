module audioControlTest


endmodule