// Test top module for ANTIC

`include "ANTIC.v"
`include "RAM.v"
`include "memoryMap.v"

module testANTIC(CPU_data);

  inout [7:0] CPU_data;

  reg reset;
  reg Fphi0;
  reg phi2;
  reg [7:0] i;      // Remember to change this accordingly
  
  wire [2:0] AN;
  wire halt_L;
  wire [15:0] address;
  wire [7:0] DB;
  wire [15:0] dlistptr;
  wire [2:0] curr_state;
  wire [7:0] data;
  wire [7:0] IR;
  wire loadIR;
  
  wire [7:0] DMACTL;
  wire [7:0] CHACTL;
  wire [7:0] HSCROL;
  wire [7:0] VSCROL;
  wire [7:0] PMBASE;
  wire [7:0] CHBASE;
  wire [7:0] WSYNC;
  wire [7:0] NMIEN;
  wire [7:0] NMIRES_NMIST_bus;
  wire [7:0] DLISTL_bus;
  wire [7:0] DLISTH_bus;
  wire [7:0] VCOUNT;
  wire [7:0] PENH;
  wire [7:0] PENV;
  wire [2:0] ANTIC_writeEn;
  
  wire [1:0] loadDLIST;
  wire [15:0] MSR;
  wire [1:0] loadMSR_both;
  
  reg [3:0] CPU_writeEn;
  reg [7:0] writeVal;
  reg write;
  
  assign CPU_data = write ? writeVal : 8'hzz;
  
  // Instantiate Modules
  memory256x256 mem(.clock(~phi2), .enable(1'b1), .we_L(1'b1), .re_L(halt_L), .address(address), .data(DB));
  
  ANTIC antic(.Fphi0(Fphi0), .LP_L(), .RW(), .rst(reset), .phi2(phi2), .DMACTL(DMACTL), .CHACTL(CHACTL),
              .HSCROL(HSCROL), .VSCROL(VSCROL), .PMBASE(PMBASE), .CHBASE(CHBASE), .WSYNC(WSYNC), .NMIEN(NMIEN), 
              .DB(DB), .NMIRES_NMIST_bus(NMIRES_NMIST_bus), .DLISTL_bus(DLISTL_bus), .DLISTH_bus(DLISTH_bus),
              .address(address), .AN(AN), .halt_L(halt_L), .NMI_L(), .RDY_L(), .REF_L(), .RNMI_L(), .phi0(), 
              .IR_out(IR), .loadIR(loadIR), .VCOUNT(VCOUNT), .PENH(PENH), .PENV(PENV), .ANTIC_writeEn(ANTIC_writeEn), 
              .printDLIST(dlistptr), .cstate(curr_state), .data(data), .MSR(MSR), .loadDLIST_both(loadDLIST), 
              .loadMSR_both(loadMSR_both));
              
  memoryMap map(.clk(phi2), .CPU_writeEn(CPU_writeEn), .ANTIC_writeEn(ANTIC_writeEn), .CPU_addr(), .VCOUNT_in(VCOUNT),
                .PENH_in(PENH), .PENV_in(PENV), .CPU_data(CPU_data), .NMIRES_NMIST_bus(NMIRES_NMIST_bus), 
                .DLISTL_bus(DLISTL_bus), .DLISTH_bus(DLISTH_bus), .DMACTL(DMACTL), .CHACTL(CHACTL),
                .HSCROL(HSCROL), .VSCROL(VSCROL), .PMBASE(PMBASE), .CHBASE(CHBASE), .WSYNC(WSYNC), .NMIEN(NMIEN));
  
  task print;
    $display("halt_L is %b, curr_state is %b, data is %h, IR is %h, loadIR is %b, AN is %b, dlistptr is %h, loadDLIST is %b, CHBASE is %h, MSR is %h, loadMSR is %b", 
             halt_L, curr_state, data, IR, loadIR, AN, dlistptr, loadDLIST, CHBASE, MSR, loadMSR_both);
  endtask
  
  initial begin
    $display("Begin ANTIC test.");
    
    // Initialize clocks
    Fphi0 = 1'b0;
    phi2 = 1'b0;
    
    // Load DLISTPTR
    CPU_writeEn = 4'd3;
    write = 1'b1;
    writeVal = 8'h00;
    
    print; @(posedge phi2); @(negedge phi2);
    CPU_writeEn = 4'd4;
    write = 1'b1;
    writeVal = 8'hA0;
    
    print; @(posedge phi2); @(negedge phi2);
    CPU_writeEn = 4'd0;
    write = 1'b0;
    
    // Reset ANTIC FSM
    reset = 1'b1;
    print; @(posedge phi2); @(negedge phi2);
    reset = 1'b0;

    // Step through display list
    for (i=8'd0; i<8'd40; i=i+8'd1) begin
      print; @(posedge phi2); print; @(negedge phi2);
    end
    
    $display("Completed ANTIC test.");
    $finish;
  end
  
  always begin
    forever #20  phi2 = ~phi2;
  end
  
  always begin
    forever #10 Fphi0 = ~Fphi0;
  end
  
endmodule